module sdl

// va_list
[typedef]
pub struct C.va_list {}
