// Copyright(C) 2025 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module sdl

//
// SDL_keycode.h
//

// Defines constants which identify keyboard keys and modifiers.
//
// Please refer to the Best Keyboard Practices document for details on what
// this information means and how best to use it.
//
// https://wiki.libsdl.org/SDL3/BestKeyboardPractices

// The SDL virtual key representation.
//
// Values of this type are used to represent keyboard keys using the current
// layout of the keyboard. These values include Unicode values representing
// the unmodified character that would be generated by pressing the key, or an
// `SDLK_*` constant for those keys that do not generate characters.
//
// A special exception is the number keys at the top of the keyboard which map
// to SDLK_0...SDLK_9 on AZERTY layouts.
//
// Keys with the `SDLK_EXTENDED_MASK` bit set do not map to a scancode or
// unicode code point.
//
// NOTE: This datatype is available since SDL 3.2.0.
pub type Keycode = u32

// Valid key modifiers (possibly OR'd together).
//
// NOTE: This datatype is available since SDL 3.2.0.
pub type Keymod = u16

pub const sdlk_extended_mask = C.SDLK_EXTENDED_MASK // (1u << 29)

pub const sdlk_scancode_mask = C.SDLK_SCANCODE_MASK // (1u << 30)

fn C.SDL_SCANCODE_TO_KEYCODE(x int) Keycode

pub fn scancode_to_keycode(scancode Scancode) Keycode {
	return C.SDL_SCANCODE_TO_KEYCODE(int(scancode))
}

pub const sdlk_unknown = C.SDLK_UNKNOWN // 0x00000000u

pub const sdlk_return = C.SDLK_RETURN // 0x0000000du

pub const sdlk_escape = C.SDLK_ESCAPE // 0x0000001bu

pub const sdlk_backspace = C.SDLK_BACKSPACE // 0x00000008u

pub const sdlk_tab = C.SDLK_TAB // 0x00000009u

pub const sdlk_space = C.SDLK_SPACE // 0x00000020u

pub const sdlk_exclaim = C.SDLK_EXCLAIM // 0x00000021u

pub const sdlk_dblapostrophe = C.SDLK_DBLAPOSTROPHE // 0x00000022u

pub const sdlk_hash = C.SDLK_HASH // 0x00000023u

pub const sdlk_dollar = C.SDLK_DOLLAR // 0x00000024u

pub const sdlk_percent = C.SDLK_PERCENT // 0x00000025u

pub const sdlk_ampersand = C.SDLK_AMPERSAND // 0x00000026u

pub const sdlk_apostrophe = C.SDLK_APOSTROPHE // 0x00000027u

pub const sdlk_leftparen = C.SDLK_LEFTPAREN // 0x00000028u

pub const sdlk_rightparen = C.SDLK_RIGHTPAREN // 0x00000029u

pub const sdlk_asterisk = C.SDLK_ASTERISK // 0x0000002au

pub const sdlk_plus = C.SDLK_PLUS // 0x0000002bu

pub const sdlk_comma = C.SDLK_COMMA // 0x0000002cu

pub const sdlk_minus = C.SDLK_MINUS // 0x0000002du

pub const sdlk_period = C.SDLK_PERIOD // 0x0000002eu

pub const sdlk_slash = C.SDLK_SLASH // 0x0000002fu

pub const sdlk_0 = C.SDLK_0 // 0x00000030u

pub const sdlk_1 = C.SDLK_1 // 0x00000031u

pub const sdlk_2 = C.SDLK_2 // 0x00000032u

pub const sdlk_3 = C.SDLK_3 // 0x00000033u

pub const sdlk_4 = C.SDLK_4 // 0x00000034u

pub const sdlk_5 = C.SDLK_5 // 0x00000035u

pub const sdlk_6 = C.SDLK_6 // 0x00000036u

pub const sdlk_7 = C.SDLK_7 // 0x00000037u

pub const sdlk_8 = C.SDLK_8 // 0x00000038u

pub const sdlk_9 = C.SDLK_9 // 0x00000039u

pub const sdlk_colon = C.SDLK_COLON // 0x0000003au

pub const sdlk_semicolon = C.SDLK_SEMICOLON // 0x0000003bu

pub const sdlk_less = C.SDLK_LESS // 0x0000003cu

pub const sdlk_equals = C.SDLK_EQUALS // 0x0000003du

pub const sdlk_greater = C.SDLK_GREATER // 0x0000003eu

pub const sdlk_question = C.SDLK_QUESTION // 0x0000003fu

pub const sdlk_at = C.SDLK_AT // 0x00000040u

pub const sdlk_leftbracket = C.SDLK_LEFTBRACKET // 0x0000005bu

pub const sdlk_backslash = C.SDLK_BACKSLASH // 0x0000005cu

pub const sdlk_rightbracket = C.SDLK_RIGHTBRACKET // 0x0000005du

pub const sdlk_caret = C.SDLK_CARET // 0x0000005eu

pub const sdlk_underscore = C.SDLK_UNDERSCORE // 0x0000005fu

pub const sdlk_grave = C.SDLK_GRAVE // 0x00000060u

pub const sdlk_a = C.SDLK_A // 0x00000061u

pub const sdlk_b = C.SDLK_B // 0x00000062u

pub const sdlk_c = C.SDLK_C // 0x00000063u

pub const sdlk_d = C.SDLK_D // 0x00000064u

pub const sdlk_e = C.SDLK_E // 0x00000065u

pub const sdlk_f = C.SDLK_F // 0x00000066u

pub const sdlk_g = C.SDLK_G // 0x00000067u

pub const sdlk_h = C.SDLK_H // 0x00000068u

pub const sdlk_i = C.SDLK_I // 0x00000069u

pub const sdlk_j = C.SDLK_J // 0x0000006au

pub const sdlk_k = C.SDLK_K // 0x0000006bu

pub const sdlk_l = C.SDLK_L // 0x0000006cu

pub const sdlk_m = C.SDLK_M // 0x0000006du

pub const sdlk_n = C.SDLK_N // 0x0000006eu

pub const sdlk_o = C.SDLK_O // 0x0000006fu

pub const sdlk_p = C.SDLK_P // 0x00000070u

pub const sdlk_q = C.SDLK_Q // 0x00000071u

pub const sdlk_r = C.SDLK_R // 0x00000072u

pub const sdlk_s = C.SDLK_S // 0x00000073u

pub const sdlk_t = C.SDLK_T // 0x00000074u

pub const sdlk_u = C.SDLK_U // 0x00000075u

pub const sdlk_v = C.SDLK_V // 0x00000076u

pub const sdlk_w = C.SDLK_W // 0x00000077u

pub const sdlk_x = C.SDLK_X // 0x00000078u

pub const sdlk_y = C.SDLK_Y // 0x00000079u

pub const sdlk_z = C.SDLK_Z // 0x0000007au

pub const sdlk_leftbrace = C.SDLK_LEFTBRACE // 0x0000007bu

pub const sdlk_pipe = C.SDLK_PIPE // 0x0000007cu

pub const sdlk_rightbrace = C.SDLK_RIGHTBRACE // 0x0000007du

pub const sdlk_tilde = C.SDLK_TILDE // 0x0000007eu

pub const sdlk_delete = C.SDLK_DELETE // 0x0000007fu

pub const sdlk_plusminus = C.SDLK_PLUSMINUS // 0x000000b1u

pub const sdlk_capslock = C.SDLK_CAPSLOCK // 0x40000039u

pub const sdlk_f1 = C.SDLK_F1 // 0x4000003au

pub const sdlk_f2 = C.SDLK_F2 // 0x4000003bu

pub const sdlk_f3 = C.SDLK_F3 // 0x4000003cu

pub const sdlk_f4 = C.SDLK_F4 // 0x4000003du

pub const sdlk_f5 = C.SDLK_F5 // 0x4000003eu

pub const sdlk_f6 = C.SDLK_F6 // 0x4000003fu

pub const sdlk_f7 = C.SDLK_F7 // 0x40000040u

pub const sdlk_f8 = C.SDLK_F8 // 0x40000041u

pub const sdlk_f9 = C.SDLK_F9 // 0x40000042u

pub const sdlk_f10 = C.SDLK_F10 // 0x40000043u

pub const sdlk_f11 = C.SDLK_F11 // 0x40000044u

pub const sdlk_f12 = C.SDLK_F12 // 0x40000045u

pub const sdlk_printscreen = C.SDLK_PRINTSCREEN // 0x40000046u

pub const sdlk_scrolllock = C.SDLK_SCROLLLOCK // 0x40000047u

pub const sdlk_pause = C.SDLK_PAUSE // 0x40000048u

pub const sdlk_insert = C.SDLK_INSERT // 0x40000049u

pub const sdlk_home = C.SDLK_HOME // 0x4000004au

pub const sdlk_pageup = C.SDLK_PAGEUP // 0x4000004bu

pub const sdlk_end = C.SDLK_END // 0x4000004du

pub const sdlk_pagedown = C.SDLK_PAGEDOWN // 0x4000004eu

pub const sdlk_right = C.SDLK_RIGHT // 0x4000004fu

pub const sdlk_left = C.SDLK_LEFT // 0x40000050u

pub const sdlk_down = C.SDLK_DOWN // 0x40000051u

pub const sdlk_up = C.SDLK_UP // 0x40000052u

pub const sdlk_numlockclear = C.SDLK_NUMLOCKCLEAR // 0x40000053u

pub const sdlk_kp_divide = C.SDLK_KP_DIVIDE // 0x40000054u

pub const sdlk_kp_multiply = C.SDLK_KP_MULTIPLY // 0x40000055u

pub const sdlk_kp_minus = C.SDLK_KP_MINUS // 0x40000056u

pub const sdlk_kp_plus = C.SDLK_KP_PLUS // 0x40000057u

pub const sdlk_kp_enter = C.SDLK_KP_ENTER // 0x40000058u

pub const sdlk_kp_1 = C.SDLK_KP_1 // 0x40000059u

pub const sdlk_kp_2 = C.SDLK_KP_2 // 0x4000005au

pub const sdlk_kp_3 = C.SDLK_KP_3 // 0x4000005bu

pub const sdlk_kp_4 = C.SDLK_KP_4 // 0x4000005cu

pub const sdlk_kp_5 = C.SDLK_KP_5 // 0x4000005du

pub const sdlk_kp_6 = C.SDLK_KP_6 // 0x4000005eu

pub const sdlk_kp_7 = C.SDLK_KP_7 // 0x4000005fu

pub const sdlk_kp_8 = C.SDLK_KP_8 // 0x40000060u

pub const sdlk_kp_9 = C.SDLK_KP_9 // 0x40000061u

pub const sdlk_kp_0 = C.SDLK_KP_0 // 0x40000062u

pub const sdlk_kp_period = C.SDLK_KP_PERIOD // 0x40000063u

pub const sdlk_application = C.SDLK_APPLICATION // 0x40000065u

pub const sdlk_power = C.SDLK_POWER // 0x40000066u

pub const sdlk_kp_equals = C.SDLK_KP_EQUALS // 0x40000067u

pub const sdlk_f13 = C.SDLK_F13 // 0x40000068u

pub const sdlk_f14 = C.SDLK_F14 // 0x40000069u

pub const sdlk_f15 = C.SDLK_F15 // 0x4000006au

pub const sdlk_f16 = C.SDLK_F16 // 0x4000006bu

pub const sdlk_f17 = C.SDLK_F17 // 0x4000006cu

pub const sdlk_f18 = C.SDLK_F18 // 0x4000006du

pub const sdlk_f19 = C.SDLK_F19 // 0x4000006eu

pub const sdlk_f20 = C.SDLK_F20 // 0x4000006fu

pub const sdlk_f21 = C.SDLK_F21 // 0x40000070u

pub const sdlk_f22 = C.SDLK_F22 // 0x40000071u

pub const sdlk_f23 = C.SDLK_F23 // 0x40000072u

pub const sdlk_f24 = C.SDLK_F24 // 0x40000073u

pub const sdlk_execute = C.SDLK_EXECUTE // 0x40000074u

pub const sdlk_help = C.SDLK_HELP // 0x40000075u

pub const sdlk_menu = C.SDLK_MENU // 0x40000076u

pub const sdlk_select = C.SDLK_SELECT // 0x40000077u

pub const sdlk_stop = C.SDLK_STOP // 0x40000078u

pub const sdlk_again = C.SDLK_AGAIN // 0x40000079u

pub const sdlk_undo = C.SDLK_UNDO // 0x4000007au

pub const sdlk_cut = C.SDLK_CUT // 0x4000007bu

pub const sdlk_copy = C.SDLK_COPY // 0x4000007cu

pub const sdlk_paste = C.SDLK_PASTE // 0x4000007du

pub const sdlk_find = C.SDLK_FIND // 0x4000007eu

pub const sdlk_mute = C.SDLK_MUTE // 0x4000007fu

pub const sdlk_volumeup = C.SDLK_VOLUMEUP // 0x40000080u

pub const sdlk_volumedown = C.SDLK_VOLUMEDOWN // 0x40000081u

pub const sdlk_kp_comma = C.SDLK_KP_COMMA // 0x40000085u

pub const sdlk_kp_equalsas400 = C.SDLK_KP_EQUALSAS400 // 0x40000086u

pub const sdlk_alterase = C.SDLK_ALTERASE // 0x40000099u

pub const sdlk_sysreq = C.SDLK_SYSREQ // 0x4000009au

pub const sdlk_cancel = C.SDLK_CANCEL // 0x4000009bu

pub const sdlk_clear = C.SDLK_CLEAR // 0x4000009cu

pub const sdlk_prior = C.SDLK_PRIOR // 0x4000009du

pub const sdlk_return2 = C.SDLK_RETURN2 // 0x4000009eu

pub const sdlk_separator = C.SDLK_SEPARATOR // 0x4000009fu

pub const sdlk_out = C.SDLK_OUT // 0x400000a0u

pub const sdlk_oper = C.SDLK_OPER // 0x400000a1u

pub const sdlk_clearagain = C.SDLK_CLEARAGAIN // 0x400000a2u

pub const sdlk_crsel = C.SDLK_CRSEL // 0x400000a3u

pub const sdlk_exsel = C.SDLK_EXSEL // 0x400000a4u

pub const sdlk_kp_00 = C.SDLK_KP_00 // 0x400000b0u

pub const sdlk_kp_000 = C.SDLK_KP_000 // 0x400000b1u

pub const sdlk_thousandsseparator = C.SDLK_THOUSANDSSEPARATOR // 0x400000b2u

pub const sdlk_decimalseparator = C.SDLK_DECIMALSEPARATOR // 0x400000b3u

pub const sdlk_currencyunit = C.SDLK_CURRENCYUNIT // 0x400000b4u

pub const sdlk_currencysubunit = C.SDLK_CURRENCYSUBUNIT // 0x400000b5u

pub const sdlk_kp_leftparen = C.SDLK_KP_LEFTPAREN // 0x400000b6u

pub const sdlk_kp_rightparen = C.SDLK_KP_RIGHTPAREN // 0x400000b7u

pub const sdlk_kp_leftbrace = C.SDLK_KP_LEFTBRACE // 0x400000b8u

pub const sdlk_kp_rightbrace = C.SDLK_KP_RIGHTBRACE // 0x400000b9u

pub const sdlk_kp_tab = C.SDLK_KP_TAB // 0x400000bau

pub const sdlk_kp_backspace = C.SDLK_KP_BACKSPACE // 0x400000bbu

pub const sdlk_kp_a = C.SDLK_KP_A // 0x400000bcu

pub const sdlk_kp_b = C.SDLK_KP_B // 0x400000bdu

pub const sdlk_kp_c = C.SDLK_KP_C // 0x400000beu

pub const sdlk_kp_d = C.SDLK_KP_D // 0x400000bfu

pub const sdlk_kp_e = C.SDLK_KP_E // 0x400000c0u

pub const sdlk_kp_f = C.SDLK_KP_F // 0x400000c1u

pub const sdlk_kp_xor = C.SDLK_KP_XOR // 0x400000c2u

pub const sdlk_kp_power = C.SDLK_KP_POWER // 0x400000c3u

pub const sdlk_kp_percent = C.SDLK_KP_PERCENT // 0x400000c4u

pub const sdlk_kp_less = C.SDLK_KP_LESS // 0x400000c5u

pub const sdlk_kp_greater = C.SDLK_KP_GREATER // 0x400000c6u

pub const sdlk_kp_ampersand = C.SDLK_KP_AMPERSAND // 0x400000c7u

pub const sdlk_kp_dblampersand = C.SDLK_KP_DBLAMPERSAND // 0x400000c8u

pub const sdlk_kp_verticalbar = C.SDLK_KP_VERTICALBAR // 0x400000c9u

pub const sdlk_kp_dblverticalbar = C.SDLK_KP_DBLVERTICALBAR // 0x400000cau

pub const sdlk_kp_colon = C.SDLK_KP_COLON // 0x400000cbu

pub const sdlk_kp_hash = C.SDLK_KP_HASH // 0x400000ccu

pub const sdlk_kp_space = C.SDLK_KP_SPACE // 0x400000cdu

pub const sdlk_kp_at = C.SDLK_KP_AT // 0x400000ceu

pub const sdlk_kp_exclam = C.SDLK_KP_EXCLAM // 0x400000cfu

pub const sdlk_kp_memstore = C.SDLK_KP_MEMSTORE // 0x400000d0u

pub const sdlk_kp_memrecall = C.SDLK_KP_MEMRECALL // 0x400000d1u

pub const sdlk_kp_memclear = C.SDLK_KP_MEMCLEAR // 0x400000d2u

pub const sdlk_kp_memadd = C.SDLK_KP_MEMADD // 0x400000d3u

pub const sdlk_kp_memsubtract = C.SDLK_KP_MEMSUBTRACT // 0x400000d4u

pub const sdlk_kp_memmultiply = C.SDLK_KP_MEMMULTIPLY // 0x400000d5u

pub const sdlk_kp_memdivide = C.SDLK_KP_MEMDIVIDE // 0x400000d6u

pub const sdlk_kp_plusminus = C.SDLK_KP_PLUSMINUS // 0x400000d7u

pub const sdlk_kp_clear = C.SDLK_KP_CLEAR // 0x400000d8u

pub const sdlk_kp_clearentry = C.SDLK_KP_CLEARENTRY // 0x400000d9u

pub const sdlk_kp_binary = C.SDLK_KP_BINARY // 0x400000dau

pub const sdlk_kp_octal = C.SDLK_KP_OCTAL // 0x400000dbu

pub const sdlk_kp_decimal = C.SDLK_KP_DECIMAL // 0x400000dcu

pub const sdlk_kp_hexadecimal = C.SDLK_KP_HEXADECIMAL // 0x400000ddu

pub const sdlk_lctrl = C.SDLK_LCTRL // 0x400000e0u

pub const sdlk_lshift = C.SDLK_LSHIFT // 0x400000e1u

pub const sdlk_lalt = C.SDLK_LALT // 0x400000e2u

pub const sdlk_lgui = C.SDLK_LGUI // 0x400000e3u

pub const sdlk_rctrl = C.SDLK_RCTRL // 0x400000e4u

pub const sdlk_rshift = C.SDLK_RSHIFT // 0x400000e5u

pub const sdlk_ralt = C.SDLK_RALT // 0x400000e6u

pub const sdlk_rgui = C.SDLK_RGUI // 0x400000e7u

pub const sdlk_mode = C.SDLK_MODE // 0x40000101u

pub const sdlk_sleep = C.SDLK_SLEEP // 0x40000102u

pub const sdlk_wake = C.SDLK_WAKE // 0x40000103u

pub const sdlk_channel_increment = C.SDLK_CHANNEL_INCREMENT // 0x40000104u

pub const sdlk_channel_decrement = C.SDLK_CHANNEL_DECREMENT // 0x40000105u

pub const sdlk_media_play = C.SDLK_MEDIA_PLAY // 0x40000106u

pub const sdlk_media_pause = C.SDLK_MEDIA_PAUSE // 0x40000107u

pub const sdlk_media_record = C.SDLK_MEDIA_RECORD // 0x40000108u

pub const sdlk_media_fast_forward = C.SDLK_MEDIA_FAST_FORWARD // 0x40000109u

pub const sdlk_media_rewind = C.SDLK_MEDIA_REWIND // 0x4000010au

pub const sdlk_media_next_track = C.SDLK_MEDIA_NEXT_TRACK // 0x4000010bu

pub const sdlk_media_previous_track = C.SDLK_MEDIA_PREVIOUS_TRACK // 0x4000010cu

pub const sdlk_media_stop = C.SDLK_MEDIA_STOP // 0x4000010du

pub const sdlk_media_eject = C.SDLK_MEDIA_EJECT // 0x4000010eu

pub const sdlk_media_play_pause = C.SDLK_MEDIA_PLAY_PAUSE // 0x4000010fu

pub const sdlk_media_select = C.SDLK_MEDIA_SELECT // 0x40000110u

pub const sdlk_ac_new = C.SDLK_AC_NEW // 0x40000111u

pub const sdlk_ac_open = C.SDLK_AC_OPEN // 0x40000112u

pub const sdlk_ac_close = C.SDLK_AC_CLOSE // 0x40000113u

pub const sdlk_ac_exit = C.SDLK_AC_EXIT // 0x40000114u

pub const sdlk_ac_save = C.SDLK_AC_SAVE // 0x40000115u

pub const sdlk_ac_print = C.SDLK_AC_PRINT // 0x40000116u

pub const sdlk_ac_properties = C.SDLK_AC_PROPERTIES // 0x40000117u

pub const sdlk_ac_search = C.SDLK_AC_SEARCH // 0x40000118u

pub const sdlk_ac_home = C.SDLK_AC_HOME // 0x40000119u

pub const sdlk_ac_back = C.SDLK_AC_BACK // 0x4000011au

pub const sdlk_ac_forward = C.SDLK_AC_FORWARD // 0x4000011bu

pub const sdlk_ac_stop = C.SDLK_AC_STOP // 0x4000011cu

pub const sdlk_ac_refresh = C.SDLK_AC_REFRESH // 0x4000011du

pub const sdlk_ac_bookmarks = C.SDLK_AC_BOOKMARKS // 0x4000011eu

pub const sdlk_softleft = C.SDLK_SOFTLEFT // 0x4000011fu

pub const sdlk_softright = C.SDLK_SOFTRIGHT // 0x40000120u

pub const sdlk_call = C.SDLK_CALL // 0x40000121u

pub const sdlk_endcall = C.SDLK_ENDCALL // 0x40000122u

pub const sdlk_left_tab = C.SDLK_LEFT_TAB // 0x20000001u

pub const sdlk_level5_shift = C.SDLK_LEVEL5_SHIFT // 0x20000002u

pub const sdlk_multi_key_compose = C.SDLK_MULTI_KEY_COMPOSE // 0x20000003u

pub const sdlk_lmeta = C.SDLK_LMETA // 0x20000004u

pub const sdlk_rmeta = C.SDLK_RMETA // 0x20000005u

pub const sdlk_lhyper = C.SDLK_LHYPER // 0x20000006u

pub const sdlk_rhyper = C.SDLK_RHYPER // 0x20000007u

pub const kmod_none = C.SDL_KMOD_NONE // 0x0000u

pub const kmod_lshift = C.SDL_KMOD_LSHIFT // 0x0001u

pub const kmod_rshift = C.SDL_KMOD_RSHIFT // 0x0002u

pub const kmod_level5 = C.SDL_KMOD_LEVEL5 // 0x0004u

pub const kmod_lctrl = C.SDL_KMOD_LCTRL // 0x0040u

pub const kmod_rctrl = C.SDL_KMOD_RCTRL // 0x0080u

pub const kmod_lalt = C.SDL_KMOD_LALT // 0x0100u

pub const kmod_ralt = C.SDL_KMOD_RALT // 0x0200u

pub const kmod_lgui = C.SDL_KMOD_LGUI // 0x0400u

pub const kmod_rgui = C.SDL_KMOD_RGUI // 0x0800u

pub const kmod_num = C.SDL_KMOD_NUM // 0x1000u

pub const kmod_caps = C.SDL_KMOD_CAPS // 0x2000u

pub const kmod_mode = C.SDL_KMOD_MODE // 0x4000u

pub const kmod_scroll = C.SDL_KMOD_SCROLL // 0x8000u

pub const kmod_ctrl = C.SDL_KMOD_CTRL // (SDL_KMOD_LCTRL | SDL_KMOD_RCTRL)

pub const kmod_shift = C.SDL_KMOD_SHIFT // (SDL_KMOD_LSHIFT | SDL_KMOD_RSHIFT)

pub const kmod_alt = C.SDL_KMOD_ALT // (SDL_KMOD_LALT | SDL_KMOD_RALT)

pub const kmod_gui = C.SDL_KMOD_GUI // (SDL_KMOD_LGUI | SDL_KMOD_RGUI)

// KeyMod is a convenience enum provided by the V wrapper to make modification key matching
// via `match` statements a bit easier.
pub enum KeyMod as u16 {
	none   = C.SDL_KMOD_NONE   // 0x0000u
	lshift = C.SDL_KMOD_LSHIFT // 0x0001u
	rshift = C.SDL_KMOD_RSHIFT // 0x0002u
	level5 = C.SDL_KMOD_LEVEL5 // 0x0004u
	lctrl  = C.SDL_KMOD_LCTRL  // 0x0040u
	rctrl  = C.SDL_KMOD_RCTRL  // 0x0080u
	lalt   = C.SDL_KMOD_LALT   // 0x0100u
	ralt   = C.SDL_KMOD_RALT   // 0x0200u
	lgui   = C.SDL_KMOD_LGUI   // 0x0400u
	rgui   = C.SDL_KMOD_RGUI   // 0x0800u
	num    = C.SDL_KMOD_NUM    // 0x1000u / Num-lock
	caps   = C.SDL_KMOD_CAPS   // 0x2000u / Caps-lock
	mode   = C.SDL_KMOD_MODE   // 0x4000u
	scroll = C.SDL_KMOD_SCROLL // 0x8000u / Scroll-lock
	ctrl   = C.SDL_KMOD_CTRL   // (SDL_KMOD_LCTRL | SDL_KMOD_RCTRL)
	shift  = C.SDL_KMOD_SHIFT  // (SDL_KMOD_LSHIFT | SDL_KMOD_RSHIFT)
	alt    = C.SDL_KMOD_ALT    // (SDL_KMOD_LALT | SDL_KMOD_RALT)
	gui    = C.SDL_KMOD_GUI    // (SDL_KMOD_LGUI | SDL_KMOD_RGUI)
}

// KeyCode is a convenience enum provided by the V wrapper to make key matching
// via `match` statements a bit easier.
pub enum KeyCode as u32 {
	unknown       = C.SDLK_UNKNOWN       // 0      / 0x00000000u
	return        = C.SDLK_RETURN        // `\r`   / 0x0000000du
	escape        = C.SDLK_ESCAPE        // `\x1B` / 0x0000001bu
	backspace     = C.SDLK_BACKSPACE     // `\b`   / 0x00000008u
	tab           = C.SDLK_TAB           // `\t`   / 0x00000009u
	space         = C.SDLK_SPACE         // ` `    / 0x00000020u
	exclaim       = C.SDLK_EXCLAIM       // `!`    / 0x00000021u
	dblapostrophe = C.SDLK_DBLAPOSTROPHE // `"`    / 0x00000022u
	hash          = C.SDLK_HASH          // `#`    / 0x00000023u
	dollar        = C.SDLK_DOLLAR        // `$`    / 0x00000024u
	percent       = C.SDLK_PERCENT       // `%`    / 0x00000025u
	ampersand     = C.SDLK_AMPERSAND     // `&`    / 0x00000026u
	apostrophe    = C.SDLK_APOSTROPHE    // `'`    / 0x00000027u

	leftparen  = C.SDLK_LEFTPAREN  // `(` / 0x00000028u
	rightparen = C.SDLK_RIGHTPAREN // `)` / 0x00000029u
	asterisk   = C.SDLK_ASTERISK   // `*` / 0x0000002au
	plus       = C.SDLK_PLUS       // `+` / 0x0000002bu
	comma      = C.SDLK_COMMA      // `'` / 0x0000002cu
	minus      = C.SDLK_MINUS      // `-` / 0x0000002du
	period     = C.SDLK_PERIOD     // `.` / 0x0000002eu
	slash      = C.SDLK_SLASH      // `/` / 0x0000002fu
	_0         = C.SDLK_0          // `0` / 0x00000030u
	_1         = C.SDLK_1          // `1` / 0x00000031u
	_2         = C.SDLK_2          // `2` / 0x00000032u
	_3         = C.SDLK_3          // `3` / 0x00000033u
	_4         = C.SDLK_4          // `4` / 0x00000034u
	_5         = C.SDLK_5          // `5` / 0x00000035u
	_6         = C.SDLK_6          // `6` / 0x00000036u
	_7         = C.SDLK_7          // `7` / 0x00000037u
	_8         = C.SDLK_8          // `8` / 0x00000038u
	_9         = C.SDLK_9          // `9` / 0x00000039u

	colon     = C.SDLK_COLON     // `:` / 0x0000003au
	semicolon = C.SDLK_SEMICOLON // `;` / 0x0000003bu
	less      = C.SDLK_LESS      // `<` / 0x0000003cu
	equals    = C.SDLK_EQUALS    // `=` / 0x0000003du
	greater   = C.SDLK_GREATER   // `>` / 0x0000003eu
	question  = C.SDLK_QUESTION  // `?` / 0x0000003fu
	at        = C.SDLK_AT        // `@` / 0x00000040u
	//
	leftbracket  = C.SDLK_LEFTBRACKET  // `[`  / 0x0000005bu
	backslash    = C.SDLK_BACKSLASH    // `\\` / 0x0000005cu
	rightbracket = C.SDLK_RIGHTBRACKET // `]`  / 0x0000005du
	caret        = C.SDLK_CARET        // `^`  / 0x0000005eu
	underscore   = C.SDLK_UNDERSCORE   // `_`  / 0x0000005fu
	grave        = C.SDLK_GRAVE        // `\`` / 0x00000060u
	a            = C.SDLK_A            // `a`  / 0x00000061u
	b            = C.SDLK_B            // `b`  / 0x00000062u
	c            = C.SDLK_C            // `c`  / 0x00000063u
	d            = C.SDLK_D            // `d`  / 0x00000064u
	e            = C.SDLK_E            // `e`  / 0x00000065u
	f            = C.SDLK_F            // `f`  / 0x00000066u
	g            = C.SDLK_G            // `g`  / 0x00000067u
	h            = C.SDLK_H            // `h`  / 0x00000068u
	i            = C.SDLK_I            // `i`  / 0x00000069u
	j            = C.SDLK_J            // `j`  / 0x0000006au
	k            = C.SDLK_K            // `k`  / 0x0000006bu
	l            = C.SDLK_L            // `l`  / 0x0000006cu
	m            = C.SDLK_M            // `m`  / 0x0000006du
	n            = C.SDLK_N            // `n`  / 0x0000006eu
	o            = C.SDLK_O            // `o`  / 0x0000006fu
	p            = C.SDLK_P            // `p`  / 0x00000070u
	q            = C.SDLK_Q            // `q`  / 0x00000071u
	r            = C.SDLK_R            // `r`  / 0x00000072u
	s            = C.SDLK_S            // `s`  / 0x00000073u
	t            = C.SDLK_T            // `t`  / 0x00000074u
	u            = C.SDLK_U            // `u`  / 0x00000075u
	v            = C.SDLK_V            // `v`  / 0x00000076u
	w            = C.SDLK_W            // `w`  / 0x00000077u
	x            = C.SDLK_X            // `x`  / 0x00000078u
	y            = C.SDLK_Y            // `y`  / 0x00000079u
	z            = C.SDLK_Z            // `z`  / 0x0000007au
	//
	leftbrace  = C.SDLK_LEFTBRACE  // `{`         / 0x0000007bu
	pipe       = C.SDLK_PIPE       // `|`         / 0x0000007cu
	rightbrace = C.SDLK_RIGHTBRACE // `}`         / 0x0000007du
	tilde      = C.SDLK_TILDE      // `~`         / 0x0000007eu
	delete     = C.SDLK_DELETE     // `DEL`       / 0x0000007fu / `\x7F`
	plusminus  = C.SDLK_PLUSMINUS  // `+-`        / 0x000000b1u
	capslock   = C.SDLK_CAPSLOCK   // `CAPS-LOCK` / 0x40000039u
	//
	f1  = C.SDLK_F1  // `F1`  / 0x4000003au
	f2  = C.SDLK_F2  // `F2`  / 0x4000003bu
	f3  = C.SDLK_F3  // `F3`  / 0x4000003cu
	f4  = C.SDLK_F4  // `F4`  / 0x4000003du
	f5  = C.SDLK_F5  // `F5`  / 0x4000003eu
	f6  = C.SDLK_F6  // `F6`  / 0x4000003fu
	f7  = C.SDLK_F7  // `F7`  / 0x40000040u
	f8  = C.SDLK_F8  // `F8`  / 0x40000041u
	f9  = C.SDLK_F9  // `F9`  / 0x40000042u
	f10 = C.SDLK_F10 // `F10` / 0x40000043u
	f11 = C.SDLK_F11 // `F11` / 0x40000044u
	f12 = C.SDLK_F12 // `F12` / 0x40000045u
	//
	printscreen = C.SDLK_PRINTSCREEN // 0x40000046u
	scrolllock  = C.SDLK_SCROLLLOCK  // 0x40000047u
	pause       = C.SDLK_PAUSE       // 0x40000048u
	insert      = C.SDLK_INSERT      // 0x40000049u
	home        = C.SDLK_HOME        // 0x4000004au
	pageup      = C.SDLK_PAGEUP      // 0x4000004bu
	end         = C.SDLK_END         // 0x4000004du
	pagedown    = C.SDLK_PAGEDOWN    // 0x4000004eu
	right       = C.SDLK_RIGHT       // 0x4000004fu
	left        = C.SDLK_LEFT        // 0x40000050u
	down        = C.SDLK_DOWN        // 0x40000051u
	up          = C.SDLK_UP          // 0x40000052u
	//
	numlockclear = C.SDLK_NUMLOCKCLEAR // 0x40000053u
	divide       = C.SDLK_KP_DIVIDE    // 0x40000054u
	kp_multiply  = C.SDLK_KP_MULTIPLY  // 0x40000055u
	kp_minus     = C.SDLK_KP_MINUS     // 0x40000056u
	kp_plus      = C.SDLK_KP_PLUS      // 0x40000057u
	kp_enter     = C.SDLK_KP_ENTER     // 0x40000058u
	kp_1         = C.SDLK_KP_1         // 0x40000059u
	kp_2         = C.SDLK_KP_2         // 0x4000005au
	kp_3         = C.SDLK_KP_3         // 0x4000005bu
	kp_4         = C.SDLK_KP_4         // 0x4000005cu
	kp_5         = C.SDLK_KP_5         // 0x4000005du
	kp_6         = C.SDLK_KP_6         // 0x4000005eu
	kp_7         = C.SDLK_KP_7         // 0x4000005fu
	kp_8         = C.SDLK_KP_8         // 0x40000060u
	kp_9         = C.SDLK_KP_9         // 0x40000061u
	kp_0         = C.SDLK_KP_0         // 0x40000062u
	kp_period    = C.SDLK_KP_PERIOD    // 0x40000063u
	//
	application = C.SDLK_APPLICATION // 0x40000065u
	power       = C.SDLK_POWER       // 0x40000066u
	kp_equals   = C.SDLK_KP_EQUALS   // 0x40000067u
	f13         = C.SDLK_F13         // 0x40000068u
	f14         = C.SDLK_F14         // 0x40000069u
	f15         = C.SDLK_F15         // 0x4000006au
	f16         = C.SDLK_F16         // 0x4000006bu
	f17         = C.SDLK_F17         // 0x4000006cu
	f18         = C.SDLK_F18         // 0x4000006du
	f19         = C.SDLK_F19         // 0x4000006eu
	f20         = C.SDLK_F20         // 0x4000006fu
	f21         = C.SDLK_F21         // 0x40000070u
	f22         = C.SDLK_F22         // 0x40000071u
	f23         = C.SDLK_F23         // 0x40000072u
	f24         = C.SDLK_F24         // 0x40000073u

	execute     = C.SDLK_EXECUTE        // 0x40000074u
	help        = C.SDLK_HELP           // 0x40000075u
	menu        = C.SDLK_MENU           // 0x40000076u
	select      = C.SDLK_SELECT         // 0x40000077u
	stop        = C.SDLK_STOP           // 0x40000078u
	again       = C.SDLK_AGAIN          // 0x40000079u
	undo        = C.SDLK_UNDO           // 0x4000007au
	cut         = C.SDLK_CUT            // 0x4000007bu
	copy        = C.SDLK_COPY           // 0x4000007cu
	paste       = C.SDLK_PASTE          // 0x4000007du
	find        = C.SDLK_FIND           // 0x4000007eu
	mute        = C.SDLK_MUTE           // 0x4000007fu
	volumeup    = C.SDLK_VOLUMEUP       // 0x40000080u
	volumedown  = C.SDLK_VOLUMEDOWN     // 0x40000081u
	kp_comma    = C.SDLK_KP_COMMA       // 0x40000085u
	equalsas400 = C.SDLK_KP_EQUALSAS400 // 0x40000086u
	//
	alterase   = C.SDLK_ALTERASE   // 0x40000099u
	sysreq     = C.SDLK_SYSREQ     // 0x4000009au
	cancel     = C.SDLK_CANCEL     // 0x4000009bu
	clear      = C.SDLK_CLEAR      // 0x4000009cu
	prior      = C.SDLK_PRIOR      // 0x4000009du
	return2    = C.SDLK_RETURN2    // 0x4000009eu
	separator  = C.SDLK_SEPARATOR  // 0x4000009fu
	out        = C.SDLK_OUT        // 0x400000a0u
	oper       = C.SDLK_OPER       // 0x400000a1u
	clearagain = C.SDLK_CLEARAGAIN // 0x400000a2u
	crsel      = C.SDLK_CRSEL      // 0x400000a3u
	exsel      = C.SDLK_EXSEL      // 0x400000a4u
	//
	kp_00              = C.SDLK_KP_00              // 0x400000b0u
	kp_000             = C.SDLK_KP_000             // 0x400000b1u
	thousandsseparator = C.SDLK_THOUSANDSSEPARATOR // 0x400000b2u
	decimalseparator   = C.SDLK_DECIMALSEPARATOR   // 0x400000b3u
	currencyunit       = C.SDLK_CURRENCYUNIT       // 0x400000b4u
	currencysubunit    = C.SDLK_CURRENCYSUBUNIT    // 0x400000b5u
	kp_leftparen       = C.SDLK_KP_LEFTPAREN       // 0x400000b6u
	kp_rightparen      = C.SDLK_KP_RIGHTPAREN      // 0x400000b7u
	kp_leftbrace       = C.SDLK_KP_LEFTBRACE       // 0x400000b8u
	kp_rightbrace      = C.SDLK_KP_RIGHTBRACE      // 0x400000b9u
	kp_tab             = C.SDLK_KP_TAB             // 0x400000bau
	kp_backspace       = C.SDLK_KP_BACKSPACE       // 0x400000bbu
	kp_a               = C.SDLK_KP_A               // 0x400000bcu
	kp_b               = C.SDLK_KP_B               // 0x400000bdu
	kp_c               = C.SDLK_KP_C               // 0x400000beu
	kp_d               = C.SDLK_KP_D               // 0x400000bfu
	kp_e               = C.SDLK_KP_E               // 0x400000c0u
	kp_f               = C.SDLK_KP_F               // 0x400000c1u
	kp_xor             = C.SDLK_KP_XOR             // 0x400000c2u
	kp_power           = C.SDLK_KP_POWER           // 0x400000c3u
	kp_percent         = C.SDLK_KP_PERCENT         // 0x400000c4u
	kp_less            = C.SDLK_KP_LESS            // 0x400000c5u
	kp_greater         = C.SDLK_KP_GREATER         // 0x400000c6u
	kp_ampersand       = C.SDLK_KP_AMPERSAND       // 0x400000c7u
	kp_dblampersand    = C.SDLK_KP_DBLAMPERSAND    // 0x400000c8u
	kp_verticalbar     = C.SDLK_KP_VERTICALBAR     // 0x400000c9u
	kp_dblverticalbar  = C.SDLK_KP_DBLVERTICALBAR  // 0x400000cau
	kp_colon           = C.SDLK_KP_COLON           // 0x400000cbu
	kp_hash            = C.SDLK_KP_HASH            // 0x400000ccu
	kp_space           = C.SDLK_KP_SPACE           // 0x400000cdu
	kp_at              = C.SDLK_KP_AT              // 0x400000ceu
	kp_exclam          = C.SDLK_KP_EXCLAM          // 0x400000cfu
	kp_memstore        = C.SDLK_KP_MEMSTORE        // 0x400000d0u
	kp_memrecall       = C.SDLK_KP_MEMRECALL       // 0x400000d1u
	kp_memclear        = C.SDLK_KP_MEMCLEAR        // 0x400000d2u
	kp_memadd          = C.SDLK_KP_MEMADD          // 0x400000d3u
	kp_memsubtract     = C.SDLK_KP_MEMSUBTRACT     // 0x400000d4u
	kp_memmultiply     = C.SDLK_KP_MEMMULTIPLY     // 0x400000d5u
	kp_memdivide       = C.SDLK_KP_MEMDIVIDE       // 0x400000d6u
	kp_plusminus       = C.SDLK_KP_PLUSMINUS       // 0x400000d7u
	kp_clear           = C.SDLK_KP_CLEAR           // 0x400000d8u
	kp_clearentry      = C.SDLK_KP_CLEARENTRY      // 0x400000d9u
	kp_binary          = C.SDLK_KP_BINARY          // 0x400000dau
	kp_octal           = C.SDLK_KP_OCTAL           // 0x400000dbu
	kp_decimal         = C.SDLK_KP_DECIMAL         // 0x400000dcu
	kp_hexadecimal     = C.SDLK_KP_HEXADECIMAL     // 0x400000ddu
	lctrl              = C.SDLK_LCTRL              // 0x400000e0u
	lshift             = C.SDLK_LSHIFT             // 0x400000e1u
	lalt               = C.SDLK_LALT               // 0x400000e2u
	lgui               = C.SDLK_LGUI               // 0x400000e3u
	rctrl              = C.SDLK_RCTRL              // 0x400000e4u
	rshift             = C.SDLK_RSHIFT             // 0x400000e5u
	ralt               = C.SDLK_RALT               // 0x400000e6u
	rgui               = C.SDLK_RGUI               // 0x400000e7u
	//
	mode  = C.SDLK_MODE  // 0x40000101u
	sleep = C.SDLK_SLEEP // 0x40000102u
	wake  = C.SDLK_WAKE  // 0x40000103u
	//
	channel_increment    = C.SDLK_CHANNEL_INCREMENT    // 0x40000104u
	channel_decrement    = C.SDLK_CHANNEL_DECREMENT    // 0x40000105u
	media_play           = C.SDLK_MEDIA_PLAY           // 0x40000106u
	media_pause          = C.SDLK_MEDIA_PAUSE          // 0x40000107u
	media_record         = C.SDLK_MEDIA_RECORD         // 0x40000108u
	media_fast_forward   = C.SDLK_MEDIA_FAST_FORWARD   // 0x40000109u
	media_rewind         = C.SDLK_MEDIA_REWIND         // 0x4000010au
	media_next_track     = C.SDLK_MEDIA_NEXT_TRACK     // 0x4000010bu
	media_previous_track = C.SDLK_MEDIA_PREVIOUS_TRACK // 0x4000010cu
	media_stop           = C.SDLK_MEDIA_STOP           // 0x4000010du
	media_eject          = C.SDLK_MEDIA_EJECT          // 0x4000010eu
	media_play_pause     = C.SDLK_MEDIA_PLAY_PAUSE     // 0x4000010fu
	media_select         = C.SDLK_MEDIA_SELECT         // 0x40000110u
	ac_new               = C.SDLK_AC_NEW               // 0x40000111u
	ac_open              = C.SDLK_AC_OPEN              // 0x40000112u
	ac_close             = C.SDLK_AC_CLOSE             // 0x40000113u
	ac_exit              = C.SDLK_AC_EXIT              // 0x40000114u
	ac_save              = C.SDLK_AC_SAVE              // 0x40000115u
	ac_print             = C.SDLK_AC_PRINT             // 0x40000116u
	ac_properties        = C.SDLK_AC_PROPERTIES        // 0x40000117u
	ac_search            = C.SDLK_AC_SEARCH            // 0x40000118u
	ac_home              = C.SDLK_AC_HOME              // 0x40000119u
	ac_back              = C.SDLK_AC_BACK              // 0x4000011au
	ac_forward           = C.SDLK_AC_FORWARD           // 0x4000011bu
	ac_stop              = C.SDLK_AC_STOP              // 0x4000011cu
	ac_refresh           = C.SDLK_AC_REFRESH           // 0x4000011du
	ac_bookmarks         = C.SDLK_AC_BOOKMARKS         // 0x4000011eu
	softleft             = C.SDLK_SOFTLEFT             // 0x4000011fu
	softright            = C.SDLK_SOFTRIGHT            // 0x40000120u
	call                 = C.SDLK_CALL                 // 0x40000121u
	endcall              = C.SDLK_ENDCALL              // 0x40000122u
	left_tab             = C.SDLK_LEFT_TAB             // 0x20000001u
	level5_shift         = C.SDLK_LEVEL5_SHIFT         // 0x20000002u
	multi_key_compose    = C.SDLK_MULTI_KEY_COMPOSE    // 0x20000003u
	lmeta                = C.SDLK_LMETA                // 0x20000004u
	rmeta                = C.SDLK_RMETA                // 0x20000005u
	lhyper               = C.SDLK_LHYPER               // 0x20000006u
	rhyper               = C.SDLK_RHYPER               // 0x20000007u
}
