// Setup this way to make emscripten builds work with `-no-skip-unused`
module sdl

//
// SDL_system.h
//
