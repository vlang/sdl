module image

#flag linux -lSDL2_image

#flag windows -I @VMODROOT/thirdparty/SDL2_image/include
#flag windows -L @VMODROOT/thirdparty/SDL2_image/lib/x64
#flag windows -lSDL2_image

#include <SDL_image.h>
