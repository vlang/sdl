// Copyright(C) 2025 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module sdl

//
// SDL_audio.h
//

// Audio functionality for the SDL library.
//
// All audio in SDL3 revolves around SDL_AudioStream. Whether you want to play
// or record audio, convert it, stream it, buffer it, or mix it, you're going
// to be passing it through an audio stream.
//
// Audio streams are quite flexible; they can accept any amount of data at a
// time, in any supported format, and output it as needed in any other format,
// even if the data format changes on either side halfway through.
//
// An app opens an audio device and binds any number of audio streams to it,
// feeding more data to the streams as available. When the device needs more
// data, it will pull it from all bound streams and mix them together for
// playback.
//
// Audio streams can also use an app-provided callback to supply data
// on-demand, which maps pretty closely to the SDL2 audio model.
//
// SDL also provides a simple .WAV loader in SDL_LoadWAV (and SDL_LoadWAV_IO
// if you aren't reading from a file) as a basic means to load sound data into
// your program.
//
// ## Logical audio devices
//
// In SDL3, opening a physical device (like a SoundBlaster 16 Pro) gives you a
// logical device ID that you can bind audio streams to. In almost all cases,
// logical devices can be used anywhere in the API that a physical device is
// normally used. However, since each device opening generates a new logical
// device, different parts of the program (say, a VoIP library, or
// text-to-speech framework, or maybe some other sort of mixer on top of SDL)
// can have their own device opens that do not interfere with each other; each
// logical device will mix its separate audio down to a single buffer, fed to
// the physical device, behind the scenes. As many logical devices as you like
// can come and go; SDL will only have to open the physical device at the OS
// level once, and will manage all the logical devices on top of it
// internally.
//
// One other benefit of logical devices: if you don't open a specific physical
// device, instead opting for the default, SDL can automatically migrate those
// logical devices to different hardware as circumstances change: a user
// plugged in headphones? The system default changed? SDL can transparently
// migrate the logical devices to the correct physical device seamlessly and
// keep playing; the app doesn't even have to know it happened if it doesn't
// want to.
//
// ## Simplified audio
//
// As a simplified model for when a single source of audio is all that's
// needed, an app can use SDL_OpenAudioDeviceStream, which is a single
// function to open an audio device, create an audio stream, bind that stream
// to the newly-opened device, and (optionally) provide a callback for
// obtaining audio data. When using this function, the primary interface is
// the SDL_AudioStream and the device handle is mostly hidden away; destroying
// a stream created through this function will also close the device, stream
// bindings cannot be changed, etc. One other quirk of this is that the device
// is started in a _paused_ state and must be explicitly resumed; this is
// partially to offer a clean migration for SDL2 apps and partially because
// the app might have to do more setup before playback begins; in the
// non-simplified form, nothing will play until a stream is bound to a device,
// so they start _unpaused_.
//
// ## Channel layouts
//
// Audio data passing through SDL is uncompressed PCM data, interleaved. One
// can provide their own decompression through an MP3, etc, decoder, but SDL
// does not provide this directly. Each interleaved channel of data is meant
// to be in a specific order.
//
// Abbreviations:
//
// - FRONT = single mono speaker
// - FL = front left speaker
// - FR = front right speaker
// - FC = front center speaker
// - BL = back left speaker
// - BR = back right speaker
// - SR = surround right speaker
// - SL = surround left speaker
// - BC = back center speaker
// - LFE = low-frequency speaker
//
// These are listed in the order they are laid out in memory, so "FL, FR"
// means "the front left speaker is laid out in memory first, then the front
// right, then it repeats for the next audio frame".
//
// - 1 channel (mono) layout: FRONT
// - 2 channels (stereo) layout: FL, FR
// - 3 channels (2.1) layout: FL, FR, LFE
// - 4 channels (quad) layout: FL, FR, BL, BR
// - 5 channels (4.1) layout: FL, FR, LFE, BL, BR
// - 6 channels (5.1) layout: FL, FR, FC, LFE, BL, BR (last two can also be
//   SL, SR)
// - 7 channels (6.1) layout: FL, FR, FC, LFE, BC, SL, SR
// - 8 channels (7.1) layout: FL, FR, FC, LFE, BL, BR, SL, SR
//
// This is the same order as DirectSound expects, but applied to all
// platforms; SDL will swizzle the channels as necessary if a platform expects
// something different.
//
// SDL_AudioStream can also be provided channel maps to change this ordering
// to whatever is necessary, in other audio processing scenarios.

// SDL Audio Device instance IDs.
//
// Zero is used to signify an invalid/null device.
//
// NOTE: This datatype is available since SDL 3.2.0.
pub type AudioDeviceID = u32

pub const audio_mask_bitsize = C.SDL_AUDIO_MASK_BITSIZE // (0xFFu)

pub const audio_mask_float = C.SDL_AUDIO_MASK_FLOAT // (1u<<8)

pub const audio_mask_big_endian = C.SDL_AUDIO_MASK_BIG_ENDIAN // (1u<<12)

pub const audio_mask_signed = C.SDL_AUDIO_MASK_SIGNED // (1u<<15)

// TODO: Non-numerical: #define SDL_DEFINE_AUDIO_FORMAT(signed, bigendian, flt, size) \

// AudioFormat is C.SDL_AudioFormat
pub enum AudioFormat {
	unknown = C.SDL_AUDIO_UNKNOWN // 0x0000u, Unspecified audio format
	_u8     = C.SDL_AUDIO_U8      // 0x0008u, Unsigned 8-bit samples
	_s8     = C.SDL_AUDIO_S8      // 0x8008u, Signed 8-bit samples
	_s16le  = C.SDL_AUDIO_S16LE   // 0x8010u, Signed 16-bit samples
	_s16be  = C.SDL_AUDIO_S16BE   // 0x9010u, As above, but big-endian byte order
	_s32le  = C.SDL_AUDIO_S32LE   // 0x8020u, 32-bit integer samples
	_s32be  = C.SDL_AUDIO_S32BE   // 0x9020u, As above, but big-endian byte order
	_f32le  = C.SDL_AUDIO_F32LE   // 0x8120u, 32-bit floating point samples
	_f32be  = C.SDL_AUDIO_F32BE   // 0x9120u, As above, but big-endian byte order
	_s16_1  = C.SDL_AUDIO_S16     // SDL_AUDIO_S16LE,
	_s32_1  = C.SDL_AUDIO_S32     // SDL_AUDIO_S32LE,
	_f32_1  = C.SDL_AUDIO_F32     // SDL_AUDIO_F32LE,
	_s16_2  = C.SDL_AUDIO_S16     // SDL_AUDIO_S16BE,
	_s32_2  = C.SDL_AUDIO_S32     // SDL_AUDIO_S32BE,
	_f32_2  = C.SDL_AUDIO_F32     // SDL_AUDIO_F32BE,
}

fn C.SDL_AUDIO_BITSIZE(x int) int
pub fn audio_bitsize(x int) int {
	return C.SDL_AUDIO_BITSIZE(x)
}

fn C.SDL_AUDIO_BYTESIZE(x int) int
pub fn audio_bytesize(x int) int {
	return C.SDL_AUDIO_BYTESIZE(x)
}

fn C.SDL_AUDIO_ISFLOAT(x int) bool
pub fn audio_isfloat(x int) bool {
	return C.SDL_AUDIO_ISFLOAT(x)
}

fn C.SDL_AUDIO_ISBIGENDIAN(x int) bool
pub fn audio_isbigendian(x int) bool {
	return C.SDL_AUDIO_ISBIGENDIAN(x)
}

fn C.SDL_AUDIO_ISLITTLEENDIAN(x int) bool
pub fn audio_islittleendian(x int) bool {
	return C.SDL_AUDIO_ISLITTLEENDIAN(x)
}

fn C.SDL_AUDIO_ISSIGNED(x int) bool
pub fn audio_issigned(x int) bool {
	return C.SDL_AUDIO_ISSIGNED(x)
}

fn C.SDL_AUDIO_ISINT(x int) bool
pub fn audio_isint(x int) bool {
	return C.SDL_AUDIO_ISINT(x)
}

fn C.SDL_AUDIO_ISUNSIGNED(x int) bool
pub fn audio_isunsigned(x int) bool {
	return C.SDL_AUDIO_ISUNSIGNED(x)
}

pub const audio_device_default_playback = C.SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK // ((SDL_AudioDeviceID) 0xFFFFFFFFu)

pub const audio_device_default_recording = C.SDL_AUDIO_DEVICE_DEFAULT_RECORDING // ((SDL_AudioDeviceID) 0xFFFFFFFEu)

@[typedef]
pub struct C.SDL_AudioSpec {
pub mut:
	format   AudioFormat // Audio data format
	channels int         // Number of channels: 1 mono, 2 stereo, etc
	freq     int         // sample rate: sample frames per second
}

pub type AudioSpec = C.SDL_AudioSpec

// TODO: Function: #define SDL_AUDIO_FRAMESIZE(x) (SDL_AUDIO_BYTESIZE((x).format) * (x).channels)

@[noinit; typedef]
pub struct C.SDL_AudioStream {
	// NOTE: Opaque type
}

pub type AudioStream = C.SDL_AudioStream

// C.SDL_GetNumAudioDrivers [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetNumAudioDrivers)
fn C.SDL_GetNumAudioDrivers() int

// get_num_audio_drivers uses this function to get the number of built-in audio drivers.
//
// This function returns a hardcoded number. This never returns a negative
// value; if there are no drivers compiled into this build of SDL, this
// function returns zero. The presence of a driver in this list does not mean
// it will function, it just means SDL is capable of interacting with that
// interface. For example, a build of SDL might have esound support, but if
// there's no esound server available, SDL's esound driver would fail if used.
//
// By default, SDL tries all drivers, in its preferred order, until one is
// found to be usable.
//
// returns the number of built-in audio drivers.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_driver (SDL_GetAudioDriver)
pub fn get_num_audio_drivers() int {
	return C.SDL_GetNumAudioDrivers()
}

// C.SDL_GetAudioDriver [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioDriver)
fn C.SDL_GetAudioDriver(index int) &char

// get_audio_driver uses this function to get the name of a built in audio driver.
//
// The list of audio drivers is given in the order that they are normally
// initialized by default; the drivers that seem more reasonable to choose
// first (as far as the SDL developers believe) are earlier in the list.
//
// The names of drivers are all simple, low-ASCII identifiers, like "alsa",
// "coreaudio" or "wasapi". These never have Unicode characters, and are not
// meant to be proper names.
//
// `index` index the index of the audio driver; the value ranges from 0 to
//              SDL_GetNumAudioDrivers() - 1.
// returns the name of the audio driver at the requested index, or NULL if an
//          invalid index was specified.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_num_audio_drivers (SDL_GetNumAudioDrivers)
pub fn get_audio_driver(index int) &char {
	return &char(C.SDL_GetAudioDriver(index))
}

// C.SDL_GetCurrentAudioDriver [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetCurrentAudioDriver)
fn C.SDL_GetCurrentAudioDriver() &char

// get_current_audio_driver gets the name of the current audio driver.
//
// The names of drivers are all simple, low-ASCII identifiers, like "alsa",
// "coreaudio" or "wasapi". These never have Unicode characters, and are not
// meant to be proper names.
//
// returns the name of the current audio driver or NULL if no driver has been
//          initialized.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn get_current_audio_driver() &char {
	return &char(C.SDL_GetCurrentAudioDriver())
}

// C.SDL_GetAudioPlaybackDevices [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioPlaybackDevices)
fn C.SDL_GetAudioPlaybackDevices(count &int) &AudioDeviceID

// get_audio_playback_devices gets a list of currently-connected audio playback devices.
//
// This returns of list of available devices that play sound, perhaps to
// speakers or headphones ("playback" devices). If you want devices that
// record audio, like a microphone ("recording" devices), use
// SDL_GetAudioRecordingDevices() instead.
//
// This only returns a list of physical devices; it will not have any device
// IDs returned by SDL_OpenAudioDevice().
//
// If this function returns NULL, to signify an error, `*count` will be set to
// zero.
//
// `count` count a pointer filled in with the number of devices returned, may
//              be NULL.
// returns a 0 terminated array of device instance IDs or NULL on error; call
//          SDL_GetError() for more information. This should be freed with
//          SDL_free() when it is no longer needed.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: open_audio_device (SDL_OpenAudioDevice)
// See also: get_audio_recording_devices (SDL_GetAudioRecordingDevices)
pub fn get_audio_playback_devices(count &int) &AudioDeviceID {
	return C.SDL_GetAudioPlaybackDevices(count)
}

// C.SDL_GetAudioRecordingDevices [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioRecordingDevices)
fn C.SDL_GetAudioRecordingDevices(count &int) &AudioDeviceID

// get_audio_recording_devices gets a list of currently-connected audio recording devices.
//
// This returns of list of available devices that record audio, like a
// microphone ("recording" devices). If you want devices that play sound,
// perhaps to speakers or headphones ("playback" devices), use
// SDL_GetAudioPlaybackDevices() instead.
//
// This only returns a list of physical devices; it will not have any device
// IDs returned by SDL_OpenAudioDevice().
//
// If this function returns NULL, to signify an error, `*count` will be set to
// zero.
//
// `count` count a pointer filled in with the number of devices returned, may
//              be NULL.
// returns a 0 terminated array of device instance IDs, or NULL on failure;
//          call SDL_GetError() for more information. This should be freed
//          with SDL_free() when it is no longer needed.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: open_audio_device (SDL_OpenAudioDevice)
// See also: get_audio_playback_devices (SDL_GetAudioPlaybackDevices)
pub fn get_audio_recording_devices(count &int) &AudioDeviceID {
	return C.SDL_GetAudioRecordingDevices(count)
}

// C.SDL_GetAudioDeviceName [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioDeviceName)
fn C.SDL_GetAudioDeviceName(devid AudioDeviceID) &char

// get_audio_device_name gets the human-readable name of a specific audio device.
//
// `devid` devid the instance ID of the device to query.
// returns the name of the audio device, or NULL on failure; call
//          SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_playback_devices (SDL_GetAudioPlaybackDevices)
// See also: get_audio_recording_devices (SDL_GetAudioRecordingDevices)
pub fn get_audio_device_name(devid AudioDeviceID) &char {
	return &char(C.SDL_GetAudioDeviceName(devid))
}

// C.SDL_GetAudioDeviceFormat [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioDeviceFormat)
fn C.SDL_GetAudioDeviceFormat(devid AudioDeviceID, spec &AudioSpec, sample_frames &int) bool

// get_audio_device_format gets the current audio format of a specific audio device.
//
// For an opened device, this will report the format the device is currently
// using. If the device isn't yet opened, this will report the device's
// preferred format (or a reasonable default if this can't be determined).
//
// You may also specify SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK or
// SDL_AUDIO_DEVICE_DEFAULT_RECORDING here, which is useful for getting a
// reasonable recommendation before opening the system-recommended default
// device.
//
// You can also use this to request the current device buffer size. This is
// specified in sample frames and represents the amount of data SDL will feed
// to the physical hardware in each chunk. This can be converted to
// milliseconds of audio with the following equation:
//
// `ms = (int) ((((Sint64) frames) * 1000) / spec.freq);`
//
// Buffer size is only important if you need low-level control over the audio
// playback timing. Most apps do not need this.
//
// `devid` devid the instance ID of the device to query.
// `spec` spec on return, will be filled with device details.
// `sample_frames` sample_frames pointer to store device buffer size, in sample frames.
//                      Can be NULL.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn get_audio_device_format(devid AudioDeviceID, spec &AudioSpec, sample_frames &int) bool {
	return C.SDL_GetAudioDeviceFormat(devid, spec, sample_frames)
}

// C.SDL_GetAudioDeviceChannelMap [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioDeviceChannelMap)
fn C.SDL_GetAudioDeviceChannelMap(devid AudioDeviceID, count &int) &int

// get_audio_device_channel_map gets the current channel map of an audio device.
//
// Channel maps are optional; most things do not need them, instead passing
// data in the [order that SDL expects](CategoryAudio#channel-layouts).
//
// Audio devices usually have no remapping applied. This is represented by
// returning NULL, and does not signify an error.
//
// `devid` devid the instance ID of the device to query.
// `count` count On output, set to number of channels in the map. Can be NULL.
// returns an array of the current channel mapping, with as many elements as
//          the current output spec's channels, or NULL if default. This
//          should be freed with SDL_free() when it is no longer needed.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_input_channel_map (SDL_SetAudioStreamInputChannelMap)
pub fn get_audio_device_channel_map(devid AudioDeviceID, count &int) &int {
	return C.SDL_GetAudioDeviceChannelMap(devid, count)
}

// C.SDL_OpenAudioDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_OpenAudioDevice)
fn C.SDL_OpenAudioDevice(devid AudioDeviceID, const_spec &AudioSpec) AudioDeviceID

// open_audio_device opens a specific audio device.
//
// You can open both playback and recording devices through this function.
// Playback devices will take data from bound audio streams, mix it, and send
// it to the hardware. Recording devices will feed any bound audio streams
// with a copy of any incoming data.
//
// An opened audio device starts out with no audio streams bound. To start
// audio playing, bind a stream and supply audio data to it. Unlike SDL2,
// there is no audio callback; you only bind audio streams and make sure they
// have data flowing into them (however, you can simulate SDL2's semantics
// fairly closely by using SDL_OpenAudioDeviceStream instead of this
// function).
//
// If you don't care about opening a specific device, pass a `devid` of either
// `SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK` or
// `SDL_AUDIO_DEVICE_DEFAULT_RECORDING`. In this case, SDL will try to pick
// the most reasonable default, and may also switch between physical devices
// seamlessly later, if the most reasonable default changes during the
// lifetime of this opened device (user changed the default in the OS's system
// preferences, the default got unplugged so the system jumped to a new
// default, the user plugged in headphones on a mobile device, etc). Unless
// you have a good reason to choose a specific device, this is probably what
// you want.
//
// You may request a specific format for the audio device, but there is no
// promise the device will honor that request for several reasons. As such,
// it's only meant to be a hint as to what data your app will provide. Audio
// streams will accept data in whatever format you specify and manage
// conversion for you as appropriate. SDL_GetAudioDeviceFormat can tell you
// the preferred format for the device before opening and the actual format
// the device is using after opening.
//
// It's legal to open the same device ID more than once; each successful open
// will generate a new logical SDL_AudioDeviceID that is managed separately
// from others on the same physical device. This allows libraries to open a
// device separately from the main app and bind its own streams without
// conflicting.
//
// It is also legal to open a device ID returned by a previous call to this
// function; doing so just creates another logical device on the same physical
// device. This may be useful for making logical groupings of audio streams.
//
// This function returns the opened device ID on success. This is a new,
// unique SDL_AudioDeviceID that represents a logical device.
//
// Some backends might offer arbitrary devices (for example, a networked audio
// protocol that can connect to an arbitrary server). For these, as a change
// from SDL2, you should open a default device ID and use an SDL hint to
// specify the target if you care, or otherwise let the backend figure out a
// reasonable default. Most backends don't offer anything like this, and often
// this would be an end user setting an environment variable for their custom
// need, and not something an application should specifically manage.
//
// When done with an audio device, possibly at the end of the app's life, one
// should call SDL_CloseAudioDevice() on the returned device id.
//
// `devid` devid the device instance id to open, or
//              SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK or
//              SDL_AUDIO_DEVICE_DEFAULT_RECORDING for the most reasonable
//              default device.
// `spec` spec the requested device configuration. Can be NULL to use
//             reasonable defaults.
// returns the device ID on success or 0 on failure; call SDL_GetError() for
//          more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: close_audio_device (SDL_CloseAudioDevice)
// See also: get_audio_device_format (SDL_GetAudioDeviceFormat)
pub fn open_audio_device(devid AudioDeviceID, const_spec &AudioSpec) AudioDeviceID {
	return C.SDL_OpenAudioDevice(devid, const_spec)
}

// C.SDL_IsAudioDevicePhysical [official documentation](https://wiki.libsdl.org/SDL3/SDL_IsAudioDevicePhysical)
fn C.SDL_IsAudioDevicePhysical(devid AudioDeviceID) bool

// is_audio_device_physical determines if an audio device is physical (instead of logical).
//
// An SDL_AudioDeviceID that represents physical hardware is a physical
// device; there is one for each piece of hardware that SDL can see. Logical
// devices are created by calling SDL_OpenAudioDevice or
// SDL_OpenAudioDeviceStream, and while each is associated with a physical
// device, there can be any number of logical devices on one physical device.
//
// For the most part, logical and physical IDs are interchangeable--if you try
// to open a logical device, SDL understands to assign that effort to the
// underlying physical device, etc. However, it might be useful to know if an
// arbitrary device ID is physical or logical. This function reports which.
//
// This function may return either true or false for invalid device IDs.
//
// `devid` devid the device ID to query.
// returns true if devid is a physical device, false if it is logical.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn is_audio_device_physical(devid AudioDeviceID) bool {
	return C.SDL_IsAudioDevicePhysical(devid)
}

// C.SDL_IsAudioDevicePlayback [official documentation](https://wiki.libsdl.org/SDL3/SDL_IsAudioDevicePlayback)
fn C.SDL_IsAudioDevicePlayback(devid AudioDeviceID) bool

// is_audio_device_playback determines if an audio device is a playback device (instead of recording).
//
// This function may return either true or false for invalid device IDs.
//
// `devid` devid the device ID to query.
// returns true if devid is a playback device, false if it is recording.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn is_audio_device_playback(devid AudioDeviceID) bool {
	return C.SDL_IsAudioDevicePlayback(devid)
}

// C.SDL_PauseAudioDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_PauseAudioDevice)
fn C.SDL_PauseAudioDevice(dev AudioDeviceID) bool

// pause_audio_device uses this function to pause audio playback on a specified device.
//
// This function pauses audio processing for a given device. Any bound audio
// streams will not progress, and no audio will be generated. Pausing one
// device does not prevent other unpaused devices from running.
//
// Unlike in SDL2, audio devices start in an _unpaused_ state, since an app
// has to bind a stream before any audio will flow. Pausing a paused device is
// a legal no-op.
//
// Pausing a device can be useful to halt all audio without unbinding all the
// audio streams. This might be useful while a game is paused, or a level is
// loading, etc.
//
// Physical devices can not be paused or unpaused, only logical devices
// created through SDL_OpenAudioDevice() can be.
//
// `dev` dev a device opened by SDL_OpenAudioDevice().
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: resume_audio_device (SDL_ResumeAudioDevice)
// See also: audio_device_paused (SDL_AudioDevicePaused)
pub fn pause_audio_device(dev AudioDeviceID) bool {
	return C.SDL_PauseAudioDevice(dev)
}

// C.SDL_ResumeAudioDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_ResumeAudioDevice)
fn C.SDL_ResumeAudioDevice(dev AudioDeviceID) bool

// resume_audio_device uses this function to unpause audio playback on a specified device.
//
// This function unpauses audio processing for a given device that has
// previously been paused with SDL_PauseAudioDevice(). Once unpaused, any
// bound audio streams will begin to progress again, and audio can be
// generated.
//
// Unlike in SDL2, audio devices start in an _unpaused_ state, since an app
// has to bind a stream before any audio will flow. Unpausing an unpaused
// device is a legal no-op.
//
// Physical devices can not be paused or unpaused, only logical devices
// created through SDL_OpenAudioDevice() can be.
//
// `dev` dev a device opened by SDL_OpenAudioDevice().
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: audio_device_paused (SDL_AudioDevicePaused)
// See also: pause_audio_device (SDL_PauseAudioDevice)
pub fn resume_audio_device(dev AudioDeviceID) bool {
	return C.SDL_ResumeAudioDevice(dev)
}

// C.SDL_AudioDevicePaused [official documentation](https://wiki.libsdl.org/SDL3/SDL_AudioDevicePaused)
fn C.SDL_AudioDevicePaused(dev AudioDeviceID) bool

// audio_device_paused uses this function to query if an audio device is paused.
//
// Unlike in SDL2, audio devices start in an _unpaused_ state, since an app
// has to bind a stream before any audio will flow.
//
// Physical devices can not be paused or unpaused, only logical devices
// created through SDL_OpenAudioDevice() can be. Physical and invalid device
// IDs will report themselves as unpaused here.
//
// `dev` dev a device opened by SDL_OpenAudioDevice().
// returns true if device is valid and paused, false otherwise.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: pause_audio_device (SDL_PauseAudioDevice)
// See also: resume_audio_device (SDL_ResumeAudioDevice)
pub fn audio_device_paused(dev AudioDeviceID) bool {
	return C.SDL_AudioDevicePaused(dev)
}

// C.SDL_GetAudioDeviceGain [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioDeviceGain)
fn C.SDL_GetAudioDeviceGain(devid AudioDeviceID) f32

// get_audio_device_gain gets the gain of an audio device.
//
// The gain of a device is its volume; a larger gain means a louder output,
// with a gain of zero being silence.
//
// Audio devices default to a gain of 1.0f (no change in output).
//
// Physical devices may not have their gain changed, only logical devices, and
// this function will always return -1.0f when used on physical devices.
//
// `devid` devid the audio device to query.
// returns the gain of the device or -1.0f on failure; call SDL_GetError()
//          for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_device_gain (SDL_SetAudioDeviceGain)
pub fn get_audio_device_gain(devid AudioDeviceID) f32 {
	return C.SDL_GetAudioDeviceGain(devid)
}

// C.SDL_SetAudioDeviceGain [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioDeviceGain)
fn C.SDL_SetAudioDeviceGain(devid AudioDeviceID, gain f32) bool

// set_audio_device_gain changes the gain of an audio device.
//
// The gain of a device is its volume; a larger gain means a louder output,
// with a gain of zero being silence.
//
// Audio devices default to a gain of 1.0f (no change in output).
//
// Physical devices may not have their gain changed, only logical devices, and
// this function will always return false when used on physical devices. While
// it might seem attractive to adjust several logical devices at once in this
// way, it would allow an app or library to interfere with another portion of
// the program's otherwise-isolated devices.
//
// This is applied, along with any per-audiostream gain, during playback to
// the hardware, and can be continuously changed to create various effects. On
// recording devices, this will adjust the gain before passing the data into
// an audiostream; that recording audiostream can then adjust its gain further
// when outputting the data elsewhere, if it likes, but that second gain is
// not applied until the data leaves the audiostream again.
//
// `devid` devid the audio device on which to change gain.
// `gain` gain the gain. 1.0f is no change, 0.0f is silence.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_device_gain (SDL_GetAudioDeviceGain)
pub fn set_audio_device_gain(devid AudioDeviceID, gain f32) bool {
	return C.SDL_SetAudioDeviceGain(devid, gain)
}

// C.SDL_CloseAudioDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_CloseAudioDevice)
fn C.SDL_CloseAudioDevice(devid AudioDeviceID)

// close_audio_device closes a previously-opened audio device.
//
// The application should close open audio devices once they are no longer
// needed.
//
// This function may block briefly while pending audio data is played by the
// hardware, so that applications don't drop the last buffer of data they
// supplied if terminating immediately afterwards.
//
// `devid` devid an audio device id previously returned by
//              SDL_OpenAudioDevice().
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: open_audio_device (SDL_OpenAudioDevice)
pub fn close_audio_device(devid AudioDeviceID) {
	C.SDL_CloseAudioDevice(devid)
}

// C.SDL_BindAudioStreams [official documentation](https://wiki.libsdl.org/SDL3/SDL_BindAudioStreams)
fn C.SDL_BindAudioStreams(devid AudioDeviceID, const_streams &&C.SDL_AudioStream, num_streams int) bool

// bind_audio_streams binds a list of audio streams to an audio device.
//
// Audio data will flow through any bound streams. For a playback device, data
// for all bound streams will be mixed together and fed to the device. For a
// recording device, a copy of recorded data will be provided to each bound
// stream.
//
// Audio streams can only be bound to an open device. This operation is
// atomic--all streams bound in the same call will start processing at the
// same time, so they can stay in sync. Also: either all streams will be bound
// or none of them will be.
//
// It is an error to bind an already-bound stream; it must be explicitly
// unbound first.
//
// Binding a stream to a device will set its output format for playback
// devices, and its input format for recording devices, so they match the
// device's settings. The caller is welcome to change the other end of the
// stream's format at any time with SDL_SetAudioStreamFormat().
//
// `devid` devid an audio device to bind a stream to.
// `streams` streams an array of audio streams to bind.
// `num_streams` num_streams number streams listed in the `streams` array.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: bind_audio_streams (SDL_BindAudioStreams)
// See also: unbind_audio_stream (SDL_UnbindAudioStream)
// See also: get_audio_stream_device (SDL_GetAudioStreamDevice)
pub fn bind_audio_streams(devid AudioDeviceID, const_streams &&C.SDL_AudioStream, num_streams int) bool {
	return C.SDL_BindAudioStreams(devid, voidptr(const_streams), num_streams)
}

// C.SDL_BindAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_BindAudioStream)
fn C.SDL_BindAudioStream(devid AudioDeviceID, stream &AudioStream) bool

// bind_audio_stream binds a single audio stream to an audio device.
//
// This is a convenience function, equivalent to calling
// `SDL_BindAudioStreams(devid, &stream, 1)`.
//
// `devid` devid an audio device to bind a stream to.
// `stream` stream an audio stream to bind to a device.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: bind_audio_streams (SDL_BindAudioStreams)
// See also: unbind_audio_stream (SDL_UnbindAudioStream)
// See also: get_audio_stream_device (SDL_GetAudioStreamDevice)
pub fn bind_audio_stream(devid AudioDeviceID, stream &AudioStream) bool {
	return C.SDL_BindAudioStream(devid, stream)
}

// C.SDL_UnbindAudioStreams [official documentation](https://wiki.libsdl.org/SDL3/SDL_UnbindAudioStreams)
fn C.SDL_UnbindAudioStreams(const_streams &&C.SDL_AudioStream, num_streams int)

// unbind_audio_streams unbinds a list of audio streams from their audio devices.
//
// The streams being unbound do not all have to be on the same device. All
// streams on the same device will be unbound atomically (data will stop
// flowing through all unbound streams on the same device at the same time).
//
// Unbinding a stream that isn't bound to a device is a legal no-op.
//
// `streams` streams an array of audio streams to unbind. Can be NULL or contain
//                NULL.
// `num_streams` num_streams number streams listed in the `streams` array.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: bind_audio_streams (SDL_BindAudioStreams)
pub fn unbind_audio_streams(const_streams &&C.SDL_AudioStream, num_streams int) {
	C.SDL_UnbindAudioStreams(voidptr(const_streams), num_streams)
}

// C.SDL_UnbindAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_UnbindAudioStream)
fn C.SDL_UnbindAudioStream(stream &AudioStream)

// unbind_audio_stream unbinds a single audio stream from its audio device.
//
// This is a convenience function, equivalent to calling
// `SDL_UnbindAudioStreams(&stream, 1)`.
//
// `stream` stream an audio stream to unbind from a device. Can be NULL.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: bind_audio_stream (SDL_BindAudioStream)
pub fn unbind_audio_stream(stream &AudioStream) {
	C.SDL_UnbindAudioStream(stream)
}

// C.SDL_GetAudioStreamDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamDevice)
fn C.SDL_GetAudioStreamDevice(stream &AudioStream) AudioDeviceID

// get_audio_stream_device querys an audio stream for its currently-bound device.
//
// This reports the audio device that an audio stream is currently bound to.
//
// If not bound, or invalid, this returns zero, which is not a valid device
// ID.
//
// `stream` stream the audio stream to query.
// returns the bound audio device, or 0 if not bound or invalid.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: bind_audio_stream (SDL_BindAudioStream)
// See also: bind_audio_streams (SDL_BindAudioStreams)
pub fn get_audio_stream_device(stream &AudioStream) AudioDeviceID {
	return C.SDL_GetAudioStreamDevice(stream)
}

// C.SDL_CreateAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_CreateAudioStream)
fn C.SDL_CreateAudioStream(const_src_spec &AudioSpec, const_dst_spec &AudioSpec) &AudioStream

// create_audio_stream creates a new audio stream.
//
// `src_spec` src_spec the format details of the input audio.
// `dst_spec` dst_spec the format details of the output audio.
// returns a new audio stream on success or NULL on failure; call
//          SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
// See also: get_audio_stream_data (SDL_GetAudioStreamData)
// See also: get_audio_stream_available (SDL_GetAudioStreamAvailable)
// See also: flush_audio_stream (SDL_FlushAudioStream)
// See also: clear_audio_stream (SDL_ClearAudioStream)
// See also: set_audio_stream_format (SDL_SetAudioStreamFormat)
// See also: destroy_audio_stream (SDL_DestroyAudioStream)
pub fn create_audio_stream(const_src_spec &AudioSpec, const_dst_spec &AudioSpec) &AudioStream {
	return C.SDL_CreateAudioStream(const_src_spec, const_dst_spec)
}

// C.SDL_GetAudioStreamProperties [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamProperties)
fn C.SDL_GetAudioStreamProperties(stream &AudioStream) PropertiesID

// get_audio_stream_properties gets the properties associated with an audio stream.
//
// `stream` stream the SDL_AudioStream to query.
// returns a valid property ID on success or 0 on failure; call
//          SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn get_audio_stream_properties(stream &AudioStream) PropertiesID {
	return C.SDL_GetAudioStreamProperties(stream)
}

// C.SDL_GetAudioStreamFormat [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamFormat)
fn C.SDL_GetAudioStreamFormat(stream &AudioStream, src_spec &AudioSpec, dst_spec &AudioSpec) bool

// get_audio_stream_format querys the current format of an audio stream.
//
// `stream` stream the SDL_AudioStream to query.
// `src_spec` src_spec where to store the input audio format; ignored if NULL.
// `dst_spec` dst_spec where to store the output audio format; ignored if NULL.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_format (SDL_SetAudioStreamFormat)
pub fn get_audio_stream_format(stream &AudioStream, src_spec &AudioSpec, dst_spec &AudioSpec) bool {
	return C.SDL_GetAudioStreamFormat(stream, src_spec, dst_spec)
}

// C.SDL_SetAudioStreamFormat [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamFormat)
fn C.SDL_SetAudioStreamFormat(stream &AudioStream, const_src_spec &AudioSpec, const_dst_spec &AudioSpec) bool

// set_audio_stream_format changes the input and output formats of an audio stream.
//
// Future calls to and SDL_GetAudioStreamAvailable and SDL_GetAudioStreamData
// will reflect the new format, and future calls to SDL_PutAudioStreamData
// must provide data in the new input formats.
//
// Data that was previously queued in the stream will still be operated on in
// the format that was current when it was added, which is to say you can put
// the end of a sound file in one format to a stream, change formats for the
// next sound file, and start putting that new data while the previous sound
// file is still queued, and everything will still play back correctly.
//
// If a stream is bound to a device, then the format of the side of the stream
// bound to a device cannot be changed (src_spec for recording devices,
// dst_spec for playback devices). Attempts to make a change to this side will
// be ignored, but this will not report an error. The other side's format can
// be changed.
//
// `stream` stream the stream the format is being changed.
// `src_spec` src_spec the new format of the audio input; if NULL, it is not
//                 changed.
// `dst_spec` dst_spec the new format of the audio output; if NULL, it is not
//                 changed.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_format (SDL_GetAudioStreamFormat)
// See also: set_audio_stream_frequency_ratio (SDL_SetAudioStreamFrequencyRatio)
pub fn set_audio_stream_format(stream &AudioStream, const_src_spec &AudioSpec, const_dst_spec &AudioSpec) bool {
	return C.SDL_SetAudioStreamFormat(stream, const_src_spec, const_dst_spec)
}

// C.SDL_GetAudioStreamFrequencyRatio [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamFrequencyRatio)
fn C.SDL_GetAudioStreamFrequencyRatio(stream &AudioStream) f32

// get_audio_stream_frequency_ratio gets the frequency ratio of an audio stream.
//
// `stream` stream the SDL_AudioStream to query.
// returns the frequency ratio of the stream or 0.0 on failure; call
//          SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_frequency_ratio (SDL_SetAudioStreamFrequencyRatio)
pub fn get_audio_stream_frequency_ratio(stream &AudioStream) f32 {
	return C.SDL_GetAudioStreamFrequencyRatio(stream)
}

// C.SDL_SetAudioStreamFrequencyRatio [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamFrequencyRatio)
fn C.SDL_SetAudioStreamFrequencyRatio(stream &AudioStream, ratio f32) bool

// set_audio_stream_frequency_ratio changes the frequency ratio of an audio stream.
//
// The frequency ratio is used to adjust the rate at which input data is
// consumed. Changing this effectively modifies the speed and pitch of the
// audio. A value greater than 1.0 will play the audio faster, and at a higher
// pitch. A value less than 1.0 will play the audio slower, and at a lower
// pitch.
//
// This is applied during SDL_GetAudioStreamData, and can be continuously
// changed to create various effects.
//
// `stream` stream the stream the frequency ratio is being changed.
// `ratio` ratio the frequency ratio. 1.0 is normal speed. Must be between 0.01
//              and 100.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_frequency_ratio (SDL_GetAudioStreamFrequencyRatio)
// See also: set_audio_stream_format (SDL_SetAudioStreamFormat)
pub fn set_audio_stream_frequency_ratio(stream &AudioStream, ratio f32) bool {
	return C.SDL_SetAudioStreamFrequencyRatio(stream, ratio)
}

// C.SDL_GetAudioStreamGain [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamGain)
fn C.SDL_GetAudioStreamGain(stream &AudioStream) f32

// get_audio_stream_gain gets the gain of an audio stream.
//
// The gain of a stream is its volume; a larger gain means a louder output,
// with a gain of zero being silence.
//
// Audio streams default to a gain of 1.0f (no change in output).
//
// `stream` stream the SDL_AudioStream to query.
// returns the gain of the stream or -1.0f on failure; call SDL_GetError()
//          for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_gain (SDL_SetAudioStreamGain)
pub fn get_audio_stream_gain(stream &AudioStream) f32 {
	return C.SDL_GetAudioStreamGain(stream)
}

// C.SDL_SetAudioStreamGain [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamGain)
fn C.SDL_SetAudioStreamGain(stream &AudioStream, gain f32) bool

// set_audio_stream_gain changes the gain of an audio stream.
//
// The gain of a stream is its volume; a larger gain means a louder output,
// with a gain of zero being silence.
//
// Audio streams default to a gain of 1.0f (no change in output).
//
// This is applied during SDL_GetAudioStreamData, and can be continuously
// changed to create various effects.
//
// `stream` stream the stream on which the gain is being changed.
// `gain` gain the gain. 1.0f is no change, 0.0f is silence.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_gain (SDL_GetAudioStreamGain)
pub fn set_audio_stream_gain(stream &AudioStream, gain f32) bool {
	return C.SDL_SetAudioStreamGain(stream, gain)
}

// C.SDL_GetAudioStreamInputChannelMap [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamInputChannelMap)
fn C.SDL_GetAudioStreamInputChannelMap(stream &AudioStream, count &int) &int

// get_audio_stream_input_channel_map gets the current input channel map of an audio stream.
//
// Channel maps are optional; most things do not need them, instead passing
// data in the [order that SDL expects](CategoryAudio#channel-layouts).
//
// Audio streams default to no remapping applied. This is represented by
// returning NULL, and does not signify an error.
//
// `stream` stream the SDL_AudioStream to query.
// `count` count On output, set to number of channels in the map. Can be NULL.
// returns an array of the current channel mapping, with as many elements as
//          the current output spec's channels, or NULL if default. This
//          should be freed with SDL_free() when it is no longer needed.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_input_channel_map (SDL_SetAudioStreamInputChannelMap)
pub fn get_audio_stream_input_channel_map(stream &AudioStream, count &int) &int {
	return C.SDL_GetAudioStreamInputChannelMap(stream, count)
}

// C.SDL_GetAudioStreamOutputChannelMap [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamOutputChannelMap)
fn C.SDL_GetAudioStreamOutputChannelMap(stream &AudioStream, count &int) &int

// get_audio_stream_output_channel_map gets the current output channel map of an audio stream.
//
// Channel maps are optional; most things do not need them, instead passing
// data in the [order that SDL expects](CategoryAudio#channel-layouts).
//
// Audio streams default to no remapping applied. This is represented by
// returning NULL, and does not signify an error.
//
// `stream` stream the SDL_AudioStream to query.
// `count` count On output, set to number of channels in the map. Can be NULL.
// returns an array of the current channel mapping, with as many elements as
//          the current output spec's channels, or NULL if default. This
//          should be freed with SDL_free() when it is no longer needed.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_input_channel_map (SDL_SetAudioStreamInputChannelMap)
pub fn get_audio_stream_output_channel_map(stream &AudioStream, count &int) &int {
	return C.SDL_GetAudioStreamOutputChannelMap(stream, count)
}

// C.SDL_SetAudioStreamInputChannelMap [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamInputChannelMap)
fn C.SDL_SetAudioStreamInputChannelMap(stream &AudioStream, const_chmap &int, count int) bool

// set_audio_stream_input_channel_map sets the current input channel map of an audio stream.
//
// Channel maps are optional; most things do not need them, instead passing
// data in the [order that SDL expects](CategoryAudio#channel-layouts).
//
// The input channel map reorders data that is added to a stream via
// SDL_PutAudioStreamData. Future calls to SDL_PutAudioStreamData must provide
// data in the new channel order.
//
// Each item in the array represents an input channel, and its value is the
// channel that it should be remapped to. To reverse a stereo signal's left
// and right values, you'd have an array of `{ 1, 0 }`. It is legal to remap
// multiple channels to the same thing, so `{ 1, 1 }` would duplicate the
// right channel to both channels of a stereo signal. An element in the
// channel map set to -1 instead of a valid channel will mute that channel,
// setting it to a silence value.
//
// You cannot change the number of channels through a channel map, just
// reorder/mute them.
//
// Data that was previously queued in the stream will still be operated on in
// the order that was current when it was added, which is to say you can put
// the end of a sound file in one order to a stream, change orders for the
// next sound file, and start putting that new data while the previous sound
// file is still queued, and everything will still play back correctly.
//
// Audio streams default to no remapping applied. Passing a NULL channel map
// is legal, and turns off remapping.
//
// SDL will copy the channel map; the caller does not have to save this array
// after this call.
//
// If `count` is not equal to the current number of channels in the audio
// stream's format, this will fail. This is a safety measure to make sure a
// race condition hasn't changed the format while this call is setting the
// channel map.
//
// Unlike attempting to change the stream's format, the input channel map on a
// stream bound to a recording device is permitted to change at any time; any
// data added to the stream from the device after this call will have the new
// mapping, but previously-added data will still have the prior mapping.
//
// `stream` stream the SDL_AudioStream to change.
// `chmap` chmap the new channel map, NULL to reset to default.
// `count` count The number of channels in the map.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running. Don't change the
//               stream's format to have a different number of channels from a
//               a different thread at the same time, though!
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_input_channel_map (SDL_SetAudioStreamInputChannelMap)
pub fn set_audio_stream_input_channel_map(stream &AudioStream, const_chmap &int, count int) bool {
	return C.SDL_SetAudioStreamInputChannelMap(stream, const_chmap, count)
}

// C.SDL_SetAudioStreamOutputChannelMap [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamOutputChannelMap)
fn C.SDL_SetAudioStreamOutputChannelMap(stream &AudioStream, const_chmap &int, count int) bool

// set_audio_stream_output_channel_map sets the current output channel map of an audio stream.
//
// Channel maps are optional; most things do not need them, instead passing
// data in the [order that SDL expects](CategoryAudio#channel-layouts).
//
// The output channel map reorders data that leaving a stream via
// SDL_GetAudioStreamData.
//
// Each item in the array represents an input channel, and its value is the
// channel that it should be remapped to. To reverse a stereo signal's left
// and right values, you'd have an array of `{ 1, 0 }`. It is legal to remap
// multiple channels to the same thing, so `{ 1, 1 }` would duplicate the
// right channel to both channels of a stereo signal. An element in the
// channel map set to -1 instead of a valid channel will mute that channel,
// setting it to a silence value.
//
// You cannot change the number of channels through a channel map, just
// reorder/mute them.
//
// The output channel map can be changed at any time, as output remapping is
// applied during SDL_GetAudioStreamData.
//
// Audio streams default to no remapping applied. Passing a NULL channel map
// is legal, and turns off remapping.
//
// SDL will copy the channel map; the caller does not have to save this array
// after this call.
//
// If `count` is not equal to the current number of channels in the audio
// stream's format, this will fail. This is a safety measure to make sure a
// race condition hasn't changed the format while this call is setting the
// channel map.
//
// Unlike attempting to change the stream's format, the output channel map on
// a stream bound to a recording device is permitted to change at any time;
// any data added to the stream after this call will have the new mapping, but
// previously-added data will still have the prior mapping. When the channel
// map doesn't match the hardware's channel layout, SDL will convert the data
// before feeding it to the device for playback.
//
// `stream` stream the SDL_AudioStream to change.
// `chmap` chmap the new channel map, NULL to reset to default.
// `count` count The number of channels in the map.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, as it holds
//               a stream-specific mutex while running. Don't change the
//               stream's format to have a different number of channels from a
//               a different thread at the same time, though!
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_input_channel_map (SDL_SetAudioStreamInputChannelMap)
pub fn set_audio_stream_output_channel_map(stream &AudioStream, const_chmap &int, count int) bool {
	return C.SDL_SetAudioStreamOutputChannelMap(stream, const_chmap, count)
}

// C.SDL_PutAudioStreamData [official documentation](https://wiki.libsdl.org/SDL3/SDL_PutAudioStreamData)
fn C.SDL_PutAudioStreamData(stream &AudioStream, const_buf voidptr, len int) bool

// put_audio_stream_data adds data to the stream.
//
// This data must match the format/channels/samplerate specified in the latest
// call to SDL_SetAudioStreamFormat, or the format specified when creating the
// stream if it hasn't been changed.
//
// Note that this call simply copies the unconverted data for later. This is
// different than SDL2, where data was converted during the Put call and the
// Get call would just dequeue the previously-converted data.
//
// `stream` stream the stream the audio data is being added to.
// `buf` buf a pointer to the audio data to add.
// `len` len the number of bytes to write to the stream.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, but if the
//               stream has a callback set, the caller might need to manage
//               extra locking.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: clear_audio_stream (SDL_ClearAudioStream)
// See also: flush_audio_stream (SDL_FlushAudioStream)
// See also: get_audio_stream_data (SDL_GetAudioStreamData)
// See also: get_audio_stream_queued (SDL_GetAudioStreamQueued)
pub fn put_audio_stream_data(stream &AudioStream, const_buf voidptr, len int) bool {
	return C.SDL_PutAudioStreamData(stream, const_buf, len)
}

// C.SDL_GetAudioStreamData [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamData)
fn C.SDL_GetAudioStreamData(stream &AudioStream, buf voidptr, len int) int

// get_audio_stream_data gets converted/resampled data from the stream.
//
// The input/output data format/channels/samplerate is specified when creating
// the stream, and can be changed after creation by calling
// SDL_SetAudioStreamFormat.
//
// Note that any conversion and resampling necessary is done during this call,
// and SDL_PutAudioStreamData simply queues unconverted data for later. This
// is different than SDL2, where that work was done while inputting new data
// to the stream and requesting the output just copied the converted data.
//
// `stream` stream the stream the audio is being requested from.
// `buf` buf a buffer to fill with audio data.
// `len` len the maximum number of bytes to fill.
// returns the number of bytes read from the stream or -1 on failure; call
//          SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread, but if the
//               stream has a callback set, the caller might need to manage
//               extra locking.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: clear_audio_stream (SDL_ClearAudioStream)
// See also: get_audio_stream_available (SDL_GetAudioStreamAvailable)
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
pub fn get_audio_stream_data(stream &AudioStream, buf voidptr, len int) int {
	return C.SDL_GetAudioStreamData(stream, buf, len)
}

// C.SDL_GetAudioStreamAvailable [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamAvailable)
fn C.SDL_GetAudioStreamAvailable(stream &AudioStream) int

// get_audio_stream_available gets the number of converted/resampled bytes available.
//
// The stream may be buffering data behind the scenes until it has enough to
// resample correctly, so this number might be lower than what you expect, or
// even be zero. Add more data or flush the stream if you need the data now.
//
// If the stream has so much data that it would overflow an int, the return
// value is clamped to a maximum value, but no queued data is lost; if there
// are gigabytes of data queued, the app might need to read some of it with
// SDL_GetAudioStreamData before this function's return value is no longer
// clamped.
//
// `stream` stream the audio stream to query.
// returns the number of converted/resampled bytes available or -1 on
//          failure; call SDL_GetError() for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_data (SDL_GetAudioStreamData)
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
pub fn get_audio_stream_available(stream &AudioStream) int {
	return C.SDL_GetAudioStreamAvailable(stream)
}

// C.SDL_GetAudioStreamQueued [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioStreamQueued)
fn C.SDL_GetAudioStreamQueued(stream &AudioStream) int

// get_audio_stream_queued gets the number of bytes currently queued.
//
// This is the number of bytes put into a stream as input, not the number that
// can be retrieved as output. Because of several details, it's not possible
// to calculate one number directly from the other. If you need to know how
// much usable data can be retrieved right now, you should use
// SDL_GetAudioStreamAvailable() and not this function.
//
// Note that audio streams can change their input format at any time, even if
// there is still data queued in a different format, so the returned byte
// count will not necessarily match the number of _sample frames_ available.
// Users of this API should be aware of format changes they make when feeding
// a stream and plan accordingly.
//
// Queued data is not converted until it is consumed by
// SDL_GetAudioStreamData, so this value should be representative of the exact
// data that was put into the stream.
//
// If the stream has so much data that it would overflow an int, the return
// value is clamped to a maximum value, but no queued data is lost; if there
// are gigabytes of data queued, the app might need to read some of it with
// SDL_GetAudioStreamData before this function's return value is no longer
// clamped.
//
// `stream` stream the audio stream to query.
// returns the number of bytes queued or -1 on failure; call SDL_GetError()
//          for more information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
// See also: clear_audio_stream (SDL_ClearAudioStream)
pub fn get_audio_stream_queued(stream &AudioStream) int {
	return C.SDL_GetAudioStreamQueued(stream)
}

// C.SDL_FlushAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_FlushAudioStream)
fn C.SDL_FlushAudioStream(stream &AudioStream) bool

// flush_audio_stream tells the stream that you're done sending data, and anything being buffered
// should be converted/resampled and made available immediately.
//
// It is legal to add more data to a stream after flushing, but there may be
// audio gaps in the output. Generally this is intended to signal the end of
// input, so the complete output becomes available.
//
// `stream` stream the audio stream to flush.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
pub fn flush_audio_stream(stream &AudioStream) bool {
	return C.SDL_FlushAudioStream(stream)
}

// C.SDL_ClearAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_ClearAudioStream)
fn C.SDL_ClearAudioStream(stream &AudioStream) bool

// clear_audio_stream clears any pending data in the stream.
//
// This drops any queued data, so there will be nothing to read from the
// stream until more is added.
//
// `stream` stream the audio stream to clear.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_available (SDL_GetAudioStreamAvailable)
// See also: get_audio_stream_data (SDL_GetAudioStreamData)
// See also: get_audio_stream_queued (SDL_GetAudioStreamQueued)
// See also: put_audio_stream_data (SDL_PutAudioStreamData)
pub fn clear_audio_stream(stream &AudioStream) bool {
	return C.SDL_ClearAudioStream(stream)
}

// C.SDL_PauseAudioStreamDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_PauseAudioStreamDevice)
fn C.SDL_PauseAudioStreamDevice(stream &AudioStream) bool

// pause_audio_stream_device uses this function to pause audio playback on the audio device associated
// with an audio stream.
//
// This function pauses audio processing for a given device. Any bound audio
// streams will not progress, and no audio will be generated. Pausing one
// device does not prevent other unpaused devices from running.
//
// Pausing a device can be useful to halt all audio without unbinding all the
// audio streams. This might be useful while a game is paused, or a level is
// loading, etc.
//
// `stream` stream the audio stream associated with the audio device to pause.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: resume_audio_stream_device (SDL_ResumeAudioStreamDevice)
pub fn pause_audio_stream_device(stream &AudioStream) bool {
	return C.SDL_PauseAudioStreamDevice(stream)
}

// C.SDL_ResumeAudioStreamDevice [official documentation](https://wiki.libsdl.org/SDL3/SDL_ResumeAudioStreamDevice)
fn C.SDL_ResumeAudioStreamDevice(stream &AudioStream) bool

// resume_audio_stream_device uses this function to unpause audio playback on the audio device associated
// with an audio stream.
//
// This function unpauses audio processing for a given device that has
// previously been paused. Once unpaused, any bound audio streams will begin
// to progress again, and audio can be generated.
//
// `stream` stream the audio stream associated with the audio device to resume.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: pause_audio_stream_device (SDL_PauseAudioStreamDevice)
pub fn resume_audio_stream_device(stream &AudioStream) bool {
	return C.SDL_ResumeAudioStreamDevice(stream)
}

// C.SDL_AudioStreamDevicePaused [official documentation](https://wiki.libsdl.org/SDL3/SDL_AudioStreamDevicePaused)
fn C.SDL_AudioStreamDevicePaused(stream &AudioStream) bool

// audio_stream_device_paused uses this function to query if an audio device associated with a stream is
// paused.
//
// Unlike in SDL2, audio devices start in an _unpaused_ state, since an app
// has to bind a stream before any audio will flow.
//
// `stream` stream the audio stream associated with the audio device to query.
// returns true if device is valid and paused, false otherwise.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: pause_audio_stream_device (SDL_PauseAudioStreamDevice)
// See also: resume_audio_stream_device (SDL_ResumeAudioStreamDevice)
pub fn audio_stream_device_paused(stream &AudioStream) bool {
	return C.SDL_AudioStreamDevicePaused(stream)
}

// C.SDL_LockAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_LockAudioStream)
fn C.SDL_LockAudioStream(stream &AudioStream) bool

// lock_audio_stream locks an audio stream for serialized access.
//
// Each SDL_AudioStream has an internal mutex it uses to protect its data
// structures from threading conflicts. This function allows an app to lock
// that mutex, which could be useful if registering callbacks on this stream.
//
// One does not need to lock a stream to use in it most cases, as the stream
// manages this lock internally. However, this lock is held during callbacks,
// which may run from arbitrary threads at any time, so if an app needs to
// protect shared data during those callbacks, locking the stream guarantees
// that the callback is not running while the lock is held.
//
// As this is just a wrapper over SDL_LockMutex for an internal lock; it has
// all the same attributes (recursive locks are allowed, etc).
//
// `stream` stream the audio stream to lock.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: unlock_audio_stream (SDL_UnlockAudioStream)
pub fn lock_audio_stream(stream &AudioStream) bool {
	return C.SDL_LockAudioStream(stream)
}

// C.SDL_UnlockAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_UnlockAudioStream)
fn C.SDL_UnlockAudioStream(stream &AudioStream) bool

// unlock_audio_stream unlocks an audio stream for serialized access.
//
// This unlocks an audio stream after a call to SDL_LockAudioStream.
//
// `stream` stream the audio stream to unlock.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) You should only call this from the same thread that
//               previously called SDL_LockAudioStream.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: lock_audio_stream (SDL_LockAudioStream)
pub fn unlock_audio_stream(stream &AudioStream) bool {
	return C.SDL_UnlockAudioStream(stream)
}

// AudioStreamCallback as callback that fires when data passes through an SDL_AudioStream.
//
// Apps can (optionally) register a callback with an audio stream that is
// called when data is added with SDL_PutAudioStreamData, or requested with
// SDL_GetAudioStreamData.
//
// Two values are offered here: one is the amount of additional data needed to
// satisfy the immediate request (which might be zero if the stream already
// has enough data queued) and the other is the total amount being requested.
// In a Get call triggering a Put callback, these values can be different. In
// a Put call triggering a Get callback, these values are always the same.
//
// Byte counts might be slightly overestimated due to buffering or resampling,
// and may change from call to call.
//
// This callback is not required to do anything. Generally this is useful for
// adding/reading data on demand, and the app will often put/get data as
// appropriate, but the system goes on with the data currently available to it
// if this callback does nothing.
//
// `stream` stream the SDL audio stream associated with this callback.
// `additional_amount` additional_amount the amount of data, in bytes, that is needed right
//                          now.
// `total_amount` total_amount the total amount of data requested, in bytes, that is
//                     requested or available.
// `userdata` userdata an opaque pointer provided by the app for their personal
//                 use.
//
// NOTE: (thread safety) This callbacks may run from any thread, so if you need to
//               protect shared data, you should use SDL_LockAudioStream to
//               serialize access; this lock will be held before your callback
//               is called, so your callback does not need to manage the lock
//               explicitly.
//
// NOTE: This datatype is available since SDL 3.2.0.
//
// See also: set_audio_stream_get_callback (SDL_SetAudioStreamGetCallback)
// See also: set_audio_stream_put_callback (SDL_SetAudioStreamPutCallback)
//
// [Official documentation](https://wiki.libsdl.org/SDL3/SDL_AudioStreamCallback)
pub type AudioStreamCallback = fn (userdata voidptr, stream &AudioStream, additional_amount int, total_amount int)

// C.SDL_SetAudioStreamGetCallback [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamGetCallback)
fn C.SDL_SetAudioStreamGetCallback(stream &AudioStream, callback AudioStreamCallback, userdata voidptr) bool

// set_audio_stream_get_callback sets a callback that runs when data is requested from an audio stream.
//
// This callback is called _before_ data is obtained from the stream, giving
// the callback the chance to add more on-demand.
//
// The callback can (optionally) call SDL_PutAudioStreamData() to add more
// audio to the stream during this call; if needed, the request that triggered
// this callback will obtain the new data immediately.
//
// The callback's `approx_request` argument is roughly how many bytes of
// _unconverted_ data (in the stream's input format) is needed by the caller,
// although this may overestimate a little for safety. This takes into account
// how much is already in the stream and only asks for any extra necessary to
// resolve the request, which means the callback may be asked for zero bytes,
// and a different amount on each call.
//
// The callback is not required to supply exact amounts; it is allowed to
// supply too much or too little or none at all. The caller will get what's
// available, up to the amount they requested, regardless of this callback's
// outcome.
//
// Clearing or flushing an audio stream does not call this callback.
//
// This function obtains the stream's lock, which means any existing callback
// (get or put) in progress will finish running before setting the new
// callback.
//
// Setting a NULL function turns off the callback.
//
// `stream` stream the audio stream to set the new callback on.
// `callback` callback the new callback function to call when data is requested
//                 from the stream.
// `userdata` userdata an opaque pointer provided to the callback for its own
//                 personal use.
// returns true on success or false on failure; call SDL_GetError() for more
//          information. This only fails if `stream` is NULL.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_put_callback (SDL_SetAudioStreamPutCallback)
pub fn set_audio_stream_get_callback(stream &AudioStream, callback AudioStreamCallback, userdata voidptr) bool {
	return C.SDL_SetAudioStreamGetCallback(stream, callback, userdata)
}

// C.SDL_SetAudioStreamPutCallback [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioStreamPutCallback)
fn C.SDL_SetAudioStreamPutCallback(stream &AudioStream, callback AudioStreamCallback, userdata voidptr) bool

// set_audio_stream_put_callback sets a callback that runs when data is added to an audio stream.
//
// This callback is called _after_ the data is added to the stream, giving the
// callback the chance to obtain it immediately.
//
// The callback can (optionally) call SDL_GetAudioStreamData() to obtain audio
// from the stream during this call.
//
// The callback's `approx_request` argument is how many bytes of _converted_
// data (in the stream's output format) was provided by the caller, although
// this may underestimate a little for safety. This value might be less than
// what is currently available in the stream, if data was already there, and
// might be less than the caller provided if the stream needs to keep a buffer
// to aid in resampling. Which means the callback may be provided with zero
// bytes, and a different amount on each call.
//
// The callback may call SDL_GetAudioStreamAvailable to see the total amount
// currently available to read from the stream, instead of the total provided
// by the current call.
//
// The callback is not required to obtain all data. It is allowed to read less
// or none at all. Anything not read now simply remains in the stream for
// later access.
//
// Clearing or flushing an audio stream does not call this callback.
//
// This function obtains the stream's lock, which means any existing callback
// (get or put) in progress will finish running before setting the new
// callback.
//
// Setting a NULL function turns off the callback.
//
// `stream` stream the audio stream to set the new callback on.
// `callback` callback the new callback function to call when data is added to the
//                 stream.
// `userdata` userdata an opaque pointer provided to the callback for its own
//                 personal use.
// returns true on success or false on failure; call SDL_GetError() for more
//          information. This only fails if `stream` is NULL.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: set_audio_stream_get_callback (SDL_SetAudioStreamGetCallback)
pub fn set_audio_stream_put_callback(stream &AudioStream, callback AudioStreamCallback, userdata voidptr) bool {
	return C.SDL_SetAudioStreamPutCallback(stream, callback, userdata)
}

// C.SDL_DestroyAudioStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_DestroyAudioStream)
fn C.SDL_DestroyAudioStream(stream &AudioStream)

// destroy_audio_stream frees an audio stream.
//
// This will release all allocated data, including any audio that is still
// queued. You do not need to manually clear the stream first.
//
// If this stream was bound to an audio device, it is unbound during this
// call. If this stream was created with SDL_OpenAudioDeviceStream, the audio
// device that was opened alongside this stream's creation will be closed,
// too.
//
// `stream` stream the audio stream to destroy.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: create_audio_stream (SDL_CreateAudioStream)
pub fn destroy_audio_stream(stream &AudioStream) {
	C.SDL_DestroyAudioStream(stream)
}

// C.SDL_OpenAudioDeviceStream [official documentation](https://wiki.libsdl.org/SDL3/SDL_OpenAudioDeviceStream)
fn C.SDL_OpenAudioDeviceStream(devid AudioDeviceID, const_spec &AudioSpec, callback AudioStreamCallback, userdata voidptr) &AudioStream

// open_audio_device_stream conveniences function for straightforward audio init for the common case.
//
// If all your app intends to do is provide a single source of PCM audio, this
// function allows you to do all your audio setup in a single call.
//
// This is also intended to be a clean means to migrate apps from SDL2.
//
// This function will open an audio device, create a stream and bind it.
// Unlike other methods of setup, the audio device will be closed when this
// stream is destroyed, so the app can treat the returned SDL_AudioStream as
// the only object needed to manage audio playback.
//
// Also unlike other functions, the audio device begins paused. This is to map
// more closely to SDL2-style behavior, since there is no extra step here to
// bind a stream to begin audio flowing. The audio device should be resumed
// with `SDL_ResumeAudioStreamDevice(stream);`
//
// This function works with both playback and recording devices.
//
// The `spec` parameter represents the app's side of the audio stream. That
// is, for recording audio, this will be the output format, and for playing
// audio, this will be the input format. If spec is NULL, the system will
// choose the format, and the app can use SDL_GetAudioStreamFormat() to obtain
// this information later.
//
// If you don't care about opening a specific audio device, you can (and
// probably _should_), use SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK for playback and
// SDL_AUDIO_DEVICE_DEFAULT_RECORDING for recording.
//
// One can optionally provide a callback function; if NULL, the app is
// expected to queue audio data for playback (or unqueue audio data if
// capturing). Otherwise, the callback will begin to fire once the device is
// unpaused.
//
// Destroying the returned stream with SDL_DestroyAudioStream will also close
// the audio device associated with this stream.
//
// `devid` devid an audio device to open, or SDL_AUDIO_DEVICE_DEFAULT_PLAYBACK
//              or SDL_AUDIO_DEVICE_DEFAULT_RECORDING.
// `spec` spec the audio stream's data format. Can be NULL.
// `callback` callback a callback where the app will provide new data for
//                 playback, or receive new data for recording. Can be NULL,
//                 in which case the app will need to call
//                 SDL_PutAudioStreamData or SDL_GetAudioStreamData as
//                 necessary.
// `userdata` userdata app-controlled pointer passed to callback. Can be NULL.
//                 Ignored if callback is NULL.
// returns an audio stream on success, ready to use, or NULL on failure; call
//          SDL_GetError() for more information. When done with this stream,
//          call SDL_DestroyAudioStream to free resources and close the
//          device.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: get_audio_stream_device (SDL_GetAudioStreamDevice)
// See also: resume_audio_stream_device (SDL_ResumeAudioStreamDevice)
pub fn open_audio_device_stream(devid AudioDeviceID, const_spec &AudioSpec, callback AudioStreamCallback, userdata voidptr) &AudioStream {
	return C.SDL_OpenAudioDeviceStream(devid, const_spec, callback, userdata)
}

// AudioPostmixCallback as callback that fires when data is about to be fed to an audio device.
//
// This is useful for accessing the final mix, perhaps for writing a
// visualizer or applying a final effect to the audio data before playback.
//
// This callback should run as quickly as possible and not block for any
// significant time, as this callback delays submission of data to the audio
// device, which can cause audio playback problems.
//
// The postmix callback _must_ be able to handle any audio data format
// specified in `spec`, which can change between callbacks if the audio device
// changed. However, this only covers frequency and channel count; data is
// always provided here in SDL_AUDIO_F32 format.
//
// The postmix callback runs _after_ logical device gain and audiostream gain
// have been applied, which is to say you can make the output data louder at
// this point than the gain settings would suggest.
//
// `userdata` userdata a pointer provided by the app through
//                 SDL_SetAudioPostmixCallback, for its own use.
// `spec` spec the current format of audio that is to be submitted to the
//             audio device.
// `buffer` buffer the buffer of audio samples to be submitted. The callback can
//               inspect and/or modify this data.
// `buflen` buflen the size of `buffer` in bytes.
//
// NOTE: (thread safety) This will run from a background thread owned by SDL. The
//               application is responsible for locking resources the callback
//               touches that need to be protected.
//
// NOTE: This datatype is available since SDL 3.2.0.
//
// See also: set_audio_postmix_callback (SDL_SetAudioPostmixCallback)
//
// [Official documentation](https://wiki.libsdl.org/SDL3/SDL_AudioPostmixCallback)
pub type AudioPostmixCallback = fn (userdata voidptr, const_spec &AudioSpec, buffer &f32, buflen int)

// C.SDL_SetAudioPostmixCallback [official documentation](https://wiki.libsdl.org/SDL3/SDL_SetAudioPostmixCallback)
fn C.SDL_SetAudioPostmixCallback(devid AudioDeviceID, callback AudioPostmixCallback, userdata voidptr) bool

// set_audio_postmix_callback sets a callback that fires when data is about to be fed to an audio device.
//
// This is useful for accessing the final mix, perhaps for writing a
// visualizer or applying a final effect to the audio data before playback.
//
// The buffer is the final mix of all bound audio streams on an opened device;
// this callback will fire regularly for any device that is both opened and
// unpaused. If there is no new data to mix, either because no streams are
// bound to the device or all the streams are empty, this callback will still
// fire with the entire buffer set to silence.
//
// This callback is allowed to make changes to the data; the contents of the
// buffer after this call is what is ultimately passed along to the hardware.
//
// The callback is always provided the data in float format (values from -1.0f
// to 1.0f), but the number of channels or sample rate may be different than
// the format the app requested when opening the device; SDL might have had to
// manage a conversion behind the scenes, or the playback might have jumped to
// new physical hardware when a system default changed, etc. These details may
// change between calls. Accordingly, the size of the buffer might change
// between calls as well.
//
// This callback can run at any time, and from any thread; if you need to
// serialize access to your app's data, you should provide and use a mutex or
// other synchronization device.
//
// All of this to say: there are specific needs this callback can fulfill, but
// it is not the simplest interface. Apps should generally provide audio in
// their preferred format through an SDL_AudioStream and let SDL handle the
// difference.
//
// This function is extremely time-sensitive; the callback should do the least
// amount of work possible and return as quickly as it can. The longer the
// callback runs, the higher the risk of audio dropouts or other problems.
//
// This function will block until the audio device is in between iterations,
// so any existing callback that might be running will finish before this
// function sets the new callback and returns.
//
// Setting a NULL callback function disables any previously-set callback.
//
// `devid` devid the ID of an opened audio device.
// `callback` callback a callback function to be called. Can be NULL.
// `userdata` userdata app-controlled pointer passed to callback. Can be NULL.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn set_audio_postmix_callback(devid AudioDeviceID, callback AudioPostmixCallback, userdata voidptr) bool {
	return C.SDL_SetAudioPostmixCallback(devid, callback, userdata)
}

// C.SDL_LoadWAV_IO [official documentation](https://wiki.libsdl.org/SDL3/SDL_LoadWAV_IO)
fn C.SDL_LoadWAV_IO(src &IOStream, closeio bool, spec &AudioSpec, audio_buf &&u8, audio_len &u32) bool

// load_wavio loads the audio data of a WAVE file into memory.
//
// Loading a WAVE file requires `src`, `spec`, `audio_buf` and `audio_len` to
// be valid pointers. The entire data portion of the file is then loaded into
// memory and decoded if necessary.
//
// Supported formats are RIFF WAVE files with the formats PCM (8, 16, 24, and
// 32 bits), IEEE Float (32 bits), Microsoft ADPCM and IMA ADPCM (4 bits), and
// A-law and mu-law (8 bits). Other formats are currently unsupported and
// cause an error.
//
// If this function succeeds, the return value is zero and the pointer to the
// audio data allocated by the function is written to `audio_buf` and its
// length in bytes to `audio_len`. The SDL_AudioSpec members `freq`,
// `channels`, and `format` are set to the values of the audio data in the
// buffer.
//
// It's necessary to use SDL_free() to free the audio data returned in
// `audio_buf` when it is no longer used.
//
// Because of the underspecification of the .WAV format, there are many
// problematic files in the wild that cause issues with strict decoders. To
// provide compatibility with these files, this decoder is lenient in regards
// to the truncation of the file, the fact chunk, and the size of the RIFF
// chunk. The hints `SDL_HINT_WAVE_RIFF_CHUNK_SIZE`,
// `SDL_HINT_WAVE_TRUNCATION`, and `SDL_HINT_WAVE_FACT_CHUNK` can be used to
// tune the behavior of the loading process.
//
// Any file that is invalid (due to truncation, corruption, or wrong values in
// the headers), too big, or unsupported causes an error. Additionally, any
// critical I/O error from the data source will terminate the loading process
// with an error. The function returns NULL on error and in all cases (with
// the exception of `src` being NULL), an appropriate error message will be
// set.
//
// It is required that the data source supports seeking.
//
// Example:
// ```c
// SDL_LoadWAV_IO(SDL_IOFromFile("sample.wav", "rb"), true, &spec, &buf, &len);
// ```
//
// Note that the SDL_LoadWAV function does this same thing for you, but in a
// less messy way:
//
// ```c
// SDL_LoadWAV("sample.wav", &spec, &buf, &len);
// ```
//
// `src` src the data source for the WAVE data.
// `closeio` closeio if true, calls SDL_CloseIO() on `src` before returning, even
//                in the case of an error.
// `spec` spec a pointer to an SDL_AudioSpec that will be set to the WAVE
//             data's format details on successful return.
// `audio_buf` audio_buf a pointer filled with the audio data, allocated by the
//                  function.
// `audio_len` audio_len a pointer filled with the length of the audio data buffer
//                  in bytes.
// returns true on success. `audio_buf` will be filled with a pointer to an
//          allocated buffer containing the audio data, and `audio_len` is
//          filled with the length of that audio buffer in bytes.
//
//          This function returns false if the .WAV file cannot be opened,
//          uses an unknown data format, or is corrupt; call SDL_GetError()
//          for more information.
//
//          When the application is done with the data returned in
//          `audio_buf`, it should call SDL_free() to dispose of it.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: free (SDL_free)
// See also: load_wav (SDL_LoadWAV)
pub fn load_wavio(src &IOStream, closeio bool, spec &AudioSpec, audio_buf &&u8, audio_len &u32) bool {
	return C.SDL_LoadWAV_IO(src, closeio, spec, audio_buf, audio_len)
}

// C.SDL_LoadWAV [official documentation](https://wiki.libsdl.org/SDL3/SDL_LoadWAV)
fn C.SDL_LoadWAV(const_path &char, spec &AudioSpec, audio_buf &&u8, audio_len &u32) bool

// load_wav loads a WAV from a file path.
//
// This is a convenience function that is effectively the same as:
//
// ```c
// SDL_LoadWAV_IO(SDL_IOFromFile(path, "rb"), true, spec, audio_buf, audio_len);
// ```
//
// `path` path the file path of the WAV file to open.
// `spec` spec a pointer to an SDL_AudioSpec that will be set to the WAVE
//             data's format details on successful return.
// `audio_buf` audio_buf a pointer filled with the audio data, allocated by the
//                  function.
// `audio_len` audio_len a pointer filled with the length of the audio data buffer
//                  in bytes.
// returns true on success. `audio_buf` will be filled with a pointer to an
//          allocated buffer containing the audio data, and `audio_len` is
//          filled with the length of that audio buffer in bytes.
//
//          This function returns false if the .WAV file cannot be opened,
//          uses an unknown data format, or is corrupt; call SDL_GetError()
//          for more information.
//
//          When the application is done with the data returned in
//          `audio_buf`, it should call SDL_free() to dispose of it.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
//
// See also: free (SDL_free)
// See also: load_wavio (SDL_LoadWAV_IO)
pub fn load_wav(const_path &char, spec &AudioSpec, audio_buf &&u8, audio_len &u32) bool {
	return C.SDL_LoadWAV(const_path, spec, audio_buf, audio_len)
}

// C.SDL_MixAudio [official documentation](https://wiki.libsdl.org/SDL3/SDL_MixAudio)
fn C.SDL_MixAudio(dst &u8, const_src &u8, format AudioFormat, len u32, volume f32) bool

// mix_audio mixs audio data in a specified format.
//
// This takes an audio buffer `src` of `len` bytes of `format` data and mixes
// it into `dst`, performing addition, volume adjustment, and overflow
// clipping. The buffer pointed to by `dst` must also be `len` bytes of
// `format` data.
//
// This is provided for convenience -- you can mix your own audio data.
//
// Do not use this function for mixing together more than two streams of
// sample data. The output from repeated application of this function may be
// distorted by clipping, because there is no accumulator with greater range
// than the input (not to mention this being an inefficient way of doing it).
//
// It is a common misconception that this function is required to write audio
// data to an output stream in an audio callback. While you can do that,
// SDL_MixAudio() is really only needed when you're mixing a single audio
// stream with a volume adjustment.
//
// `dst` dst the destination for the mixed audio.
// `src` src the source audio buffer to be mixed.
// `format` format the SDL_AudioFormat structure representing the desired audio
//               format.
// `len` len the length of the audio buffer in bytes.
// `volume` volume ranges from 0.0 - 1.0, and should be set to 1.0 for full
//               audio volume.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn mix_audio(dst &u8, const_src &u8, format AudioFormat, len u32, volume f32) bool {
	return C.SDL_MixAudio(dst, const_src, format, len, volume)
}

// C.SDL_ConvertAudioSamples [official documentation](https://wiki.libsdl.org/SDL3/SDL_ConvertAudioSamples)
fn C.SDL_ConvertAudioSamples(const_src_spec &AudioSpec, const_src_data &u8, src_len int, const_dst_spec &AudioSpec, dst_data &&u8, dst_len &int) bool

// convert_audio_samples converts some audio data of one format to another format.
//
// Please note that this function is for convenience, but should not be used
// to resample audio in blocks, as it will introduce audio artifacts on the
// boundaries. You should only use this function if you are converting audio
// data in its entirety in one call. If you want to convert audio in smaller
// chunks, use an SDL_AudioStream, which is designed for this situation.
//
// Internally, this function creates and destroys an SDL_AudioStream on each
// use, so it's also less efficient than using one directly, if you need to
// convert multiple times.
//
// `src_spec` src_spec the format details of the input audio.
// `src_data` src_data the audio data to be converted.
// `src_len` src_len the len of src_data.
// `dst_spec` dst_spec the format details of the output audio.
// `dst_data` dst_data will be filled with a pointer to converted audio data,
//                 which should be freed with SDL_free(). On error, it will be
//                 NULL.
// `dst_len` dst_len will be filled with the len of dst_data.
// returns true on success or false on failure; call SDL_GetError() for more
//          information.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn convert_audio_samples(const_src_spec &AudioSpec, const_src_data &u8, src_len int, const_dst_spec &AudioSpec, dst_data &&u8, dst_len &int) bool {
	return C.SDL_ConvertAudioSamples(const_src_spec, const_src_data, src_len, const_dst_spec,
		dst_data, dst_len)
}

// C.SDL_GetAudioFormatName [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetAudioFormatName)
fn C.SDL_GetAudioFormatName(format AudioFormat) &char

// get_audio_format_name gets the human readable name of an audio format.
//
// `format` format the audio format to query.
// returns the human readable name of the specified audio format or
//          "SDL_AUDIO_UNKNOWN" if the format isn't recognized.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn get_audio_format_name(format AudioFormat) &char {
	return &char(C.SDL_GetAudioFormatName(format))
}

// C.SDL_GetSilenceValueForFormat [official documentation](https://wiki.libsdl.org/SDL3/SDL_GetSilenceValueForFormat)
fn C.SDL_GetSilenceValueForFormat(format AudioFormat) int

// get_silence_value_for_format gets the appropriate memset value for silencing an audio format.
//
// The value returned by this function can be used as the second argument to
// memset (or SDL_memset) to set an audio buffer in a specific format to
// silence.
//
// `format` format the audio data format to query.
// returns a byte value that can be passed to memset.
//
// NOTE: (thread safety) It is safe to call this function from any thread.
//
// NOTE: This function is available since SDL 3.2.0.
pub fn get_silence_value_for_format(format AudioFormat) int {
	return C.SDL_GetSilenceValueForFormat(format)
}
